* NGSPICE file created from mux4to1_parax.ext - technology: sky130A

.subckt mux4to1_parax A2 A4 A1 A3 Z select1 VDD select0 nselect2 VSS
X0 VSS.t31 mux4onehot_0.x2.GN1.t2 mux4onehot_0.x2.GP1.t2 VSS.t30 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VDD.t27 mux4onehot_0.x1.nSEL0 a_617_3403# VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 Z.t13 mux4onehot_0.x2.GN3 A3.t2 VSS.t53 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X3 VDD.t36 mux4onehot_0.x2.GN2 mux4onehot_0.x2.GP2.t3 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_643_4499# select1.t0 VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X5 VSS.t4 VDD.t71 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X6 A4.t2 mux4onehot_0.x2.GP4.t4 Z.t1 VDD.t21 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X7 VDD.t23 mux4onehot_0.x2.GN4.t2 mux4onehot_0.x2.GP4.t2 VDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X8 mux4onehot_0.x2.GP3 mux4onehot_0.x2.GN3 VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 mux4onehot_0.x2.GP2.t2 mux4onehot_0.x2.GN2 VDD.t34 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X10 a_617_3403# mux4onehot_0.x1.nSEL1 VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X11 VDD.t14 VSS.t68 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X12 a_617_3403# mux4onehot_0.x1.nSEL0 a_671_3541# VSS.t19 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 A3.t0 mux4onehot_0.x2.GP3 Z.t11 VDD.t51 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X14 VDD.t48 a_617_4547# a_617_4371# VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X15 nselect2.t1 mux4onehot_0.select2 VSS.t47 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VSS.t24 select0.t0 mux4onehot_0.x1.nSEL0 VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_617_4547# select0.t1 VDD.t25 VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X18 VDD.t46 a_617_4371# mux4onehot_0.x2.GN3 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X19 a_671_3541# mux4onehot_0.x1.nSEL1 VSS.t52 VSS.t51 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X20 A4.t1 mux4onehot_0.x2.GP4.t5 Z.t2 VDD.t21 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X21 a_617_3819# a_617_3995# a_643_3947# VSS.t43 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X22 VDD.t38 a_617_3819# mux4onehot_0.x2.GN2 VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X23 mux4onehot_0.x1.nSEL0 select0.t2 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X24 nselect2.t3 mux4onehot_0.select2 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X25 VDD.t11 VSS.t69 VDD.t10 VDD.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X26 VSS.t57 mux4onehot_0.x2.GN3 mux4onehot_0.x2.GP3 VSS.t56 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 VSS.t1 select1.t1 a_617_3995# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X28 VDD.t68 select0.t3 mux4onehot_0.x1.nSEL0 VDD.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X29 mux4onehot_0.x2.GP1.t3 mux4onehot_0.x2.GN1.t3 VSS.t29 VSS.t28 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X30 VSS.t49 a_617_4371# mux4onehot_0.x2.GN3 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X31 mux4onehot_0.x1.nSEL0 select0.t4 VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 Z.t8 mux4onehot_0.x2.GN2 A2.t1 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X33 VSS.t42 a_617_3819# mux4onehot_0.x2.GN2 VSS.t41 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X34 mux4onehot_0.x2.GP4.t3 mux4onehot_0.x2.GN4.t3 VDD.t60 VDD.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 a_643_3947# select0.t5 VSS.t18 VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X36 VDD.t62 a_617_5059# mux4onehot_0.x2.GN4.t1 VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X37 VDD.t32 mux4onehot_0.x2.GN1.t4 mux4onehot_0.x2.GP1.t0 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X38 A1.t1 mux4onehot_0.x2.GP1.t4 Z.t4 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X39 a_617_3819# select0.t6 VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X40 Z.t6 mux4onehot_0.x2.GN1.t5 A1.t3 VSS.t27 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X41 Z.t7 mux4onehot_0.x2.GN2 A2.t0 VSS.t39 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X42 VSS.t26 select1.t2 mux4onehot_0.x1.nSEL1 VSS.t25 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X43 VSS.t61 a_617_5059# mux4onehot_0.x2.GN4.t0 VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X44 A2.t3 mux4onehot_0.x2.GP2.t4 Z.t14 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X45 VSS.t38 mux4onehot_0.x2.GN2 mux4onehot_0.x2.GP2.t1 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X46 Z.t9 mux4onehot_0.x2.GN4.t4 A4.t0 VSS.t40 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X47 VSS.t9 VDD.t72 VSS.t8 VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X48 VDD.t16 select1.t3 mux4onehot_0.x1.nSEL1 VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X49 mux4onehot_0.x1.nSEL1 select1.t4 VSS.t63 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X50 VSS.t16 mux4onehot_0.x2.GN4.t5 mux4onehot_0.x2.GP4.t1 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X51 mux4onehot_0.x2.GP3 mux4onehot_0.x2.GN3 VSS.t55 VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X52 mux4onehot_0.x2.GP2.t0 mux4onehot_0.x2.GN2 VSS.t36 VSS.t35 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X53 VDD.t8 VSS.t70 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X54 VSS.t13 select0.t7 a_617_4547# VSS.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X55 a_617_4371# a_617_4547# a_643_4499# VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X56 VDD.t64 select1.t5 a_617_5059# VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X57 mux4onehot_0.x1.nSEL1 select1.t6 VDD.t70 VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X58 VDD.t52 mux4onehot_0.x2.GN3 mux4onehot_0.x2.GP3 VDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X59 mux4onehot_0.x2.GP1.t1 mux4onehot_0.x2.GN1.t6 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X60 A3.t1 mux4onehot_0.x2.GP3 Z.t10 VDD.t51 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X61 a_617_5059# select0.t8 VDD.t66 VDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X62 VSS.t22 VDD.t73 VSS.t21 VSS.t20 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X63 VDD.t56 a_617_3403# mux4onehot_0.x2.GN1.t1 VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X64 VDD.t5 VSS.t71 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X65 Z.t15 mux4onehot_0.x2.GN4.t6 A4.t3 VSS.t40 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X66 a_617_5059# select1.t7 a_671_5197# VSS.t14 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X67 VSS.t45 mux4onehot_0.select2 nselect2.t0 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X68 a_617_3995# select1.t8 VDD.t58 VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X69 VDD.t40 a_617_3995# a_617_3819# VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X70 a_671_5197# select0.t9 VSS.t65 VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X71 a_617_4371# select1.t9 VDD.t2 VDD.t1 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X72 VSS.t59 a_617_3403# mux4onehot_0.x2.GN1.t0 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X73 Z.t5 mux4onehot_0.x2.GN1.t7 A1.t2 VSS.t27 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X74 A1.t0 mux4onehot_0.x2.GP1.t5 Z.t3 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X75 VDD.t42 mux4onehot_0.select2 nselect2.t2 VDD.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X76 VSS.t34 VDD.t74 VSS.t33 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X77 A2.t2 mux4onehot_0.x2.GP2.t5 Z.t0 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X78 Z.t12 mux4onehot_0.x2.GN3 A3.t3 VSS.t53 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X79 mux4onehot_0.x2.GP4.t0 mux4onehot_0.x2.GN4.t7 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 mux4onehot_0.x2.GN1.n1 mux4onehot_0.x2.GN1.t5 377.486
R1 mux4onehot_0.x2.GN1.n1 mux4onehot_0.x2.GN1.t7 374.202
R2 mux4onehot_0.x2.GN1.n7 mux4onehot_0.x2.GN1.t1 339.418
R3 mux4onehot_0.x2.GN1.n0 mux4onehot_0.x2.GN1.t0 274.06
R4 mux4onehot_0.x2.GN1.n4 mux4onehot_0.x2.GN1.t6 212.081
R5 mux4onehot_0.x2.GN1.n3 mux4onehot_0.x2.GN1.t4 212.081
R6 mux4onehot_0.x2.GN1.n5 mux4onehot_0.x2.GN1.n4 182.673
R7 mux4onehot_0.x2.GN1.n4 mux4onehot_0.x2.GN1.t3 139.78
R8 mux4onehot_0.x2.GN1.n3 mux4onehot_0.x2.GN1.t2 139.78
R9 mux4onehot_0.x2.GN1.n4 mux4onehot_0.x2.GN1.n3 61.346
R10 mux4onehot_0.x2.GN1 mux4onehot_0.x2.GN1.n5 15.8606
R11 mux4onehot_0.x2.GN1 mux4onehot_0.x2.GN1.n6 13.8044
R12 mux4onehot_0.x2.GN1.n2 mux4onehot_0.x2.GN1 11.6184
R13 mux4onehot_0.x2.GN1 mux4onehot_0.x2.GN1.n0 11.0989
R14 mux4onehot_0.x2.GN1 mux4onehot_0.x2.GN1.n2 10.8756
R15 mux4onehot_0.x2.GN1.n6 mux4onehot_0.x2.GN1 8.1246
R16 mux4onehot_0.x2.GN1.n8 mux4onehot_0.x2.GN1 6.6565
R17 mux4onehot_0.x2.GN1.n5 mux4onehot_0.x2.GN1 6.4005
R18 mux4onehot_0.x2.GN1.n0 mux4onehot_0.x2.GN1 6.1445
R19 mux4onehot_0.x2.GN1.n2 mux4onehot_0.x2.GN1 4.55738
R20 mux4onehot_0.x2.GN1.n8 mux4onehot_0.x2.GN1.n7 4.0914
R21 mux4onehot_0.x2.GN1 mux4onehot_0.x2.GN1.n8 3.61789
R22 mux4onehot_0.x2.GN1.n6 mux4onehot_0.x2.GN1 3.26325
R23 mux4onehot_0.x2.GN1.n0 mux4onehot_0.x2.GN1 2.86947
R24 mux4onehot_0.x2.GN1 mux4onehot_0.x2.GN1.n1 2.04102
R25 mux4onehot_0.x2.GN1.n7 mux4onehot_0.x2.GN1 1.74382
R26 mux4onehot_0.x2.GP1.n4 mux4onehot_0.x2.GP1.t5 450.938
R27 mux4onehot_0.x2.GP1.n4 mux4onehot_0.x2.GP1.t4 445.666
R28 mux4onehot_0.x2.GP1.n5 mux4onehot_0.x2.GP1.n3 195.832
R29 mux4onehot_0.x2.GP1.n1 mux4onehot_0.x2.GP1.n0 101.49
R30 mux4onehot_0.x2.GP1.n3 mux4onehot_0.x2.GP1.t0 26.5955
R31 mux4onehot_0.x2.GP1.n3 mux4onehot_0.x2.GP1.t1 26.5955
R32 mux4onehot_0.x2.GP1.n0 mux4onehot_0.x2.GP1.t2 24.9236
R33 mux4onehot_0.x2.GP1.n0 mux4onehot_0.x2.GP1.t3 24.9236
R34 mux4onehot_0.x2.GP1.n5 mux4onehot_0.x1.gpo0 11.8923
R35 mux4onehot_0.x1.gpo0 mux4onehot_0.x2.x1.GP 11.5413
R36 mux4onehot_0.x2.GP1.n2 mux4onehot_0.x1.x11.Y 10.7525
R37 mux4onehot_0.x1.x11.Y mux4onehot_0.x2.GP1.n5 8.09215
R38 mux4onehot_0.x2.GP1.n2 mux4onehot_0.x1.x11.Y 6.6565
R39 mux4onehot_0.x1.x11.Y mux4onehot_0.x2.GP1.n2 5.04292
R40 mux4onehot_0.x2.x1.GP mux4onehot_0.x2.GP1.n4 2.90754
R41 mux4onehot_0.x1.x11.Y mux4onehot_0.x2.GP1.n1 2.5605
R42 mux4onehot_0.x2.GP1.n1 mux4onehot_0.x1.x11.Y 1.93989
R43 VSS.n145 VSS.n22 545087
R44 VSS.n40 VSS 11981.2
R45 VSS.n147 VSS.n16 11744.7
R46 VSS.n147 VSS.n17 11744.7
R47 VSS.n151 VSS.n17 11744.7
R48 VSS.n151 VSS.n16 11744.7
R49 VSS.n158 VSS.n10 11744.7
R50 VSS.n154 VSS.n10 11744.7
R51 VSS.n158 VSS.n11 11744.7
R52 VSS.n154 VSS.n11 11744.7
R53 VSS.n167 VSS.n160 11744.7
R54 VSS.n171 VSS.n160 11744.7
R55 VSS.n167 VSS.n161 11744.7
R56 VSS.n171 VSS.n161 11744.7
R57 VSS.n179 VSS.n6 11744.7
R58 VSS.n179 VSS.n7 11744.7
R59 VSS.n178 VSS.n6 11744.7
R60 VSS.n178 VSS.n7 11744.7
R61 VSS.n166 VSS.n8 6117.99
R62 VSS.n153 VSS.n152 6083.44
R63 VSS.n172 VSS.n159 6028.93
R64 VSS.n173 VSS.n9 5416.06
R65 VSS.n174 VSS.n173 5357.62
R66 VSS.n40 VSS.n9 3878.48
R67 VSS.n146 VSS.n145 2026.31
R68 VSS.t12 VSS 1289.66
R69 VSS.n107 VSS.n41 1198.25
R70 VSS.n144 VSS.n143 1198.25
R71 VSS.n133 VSS.n29 1194.5
R72 VSS.n94 VSS.n93 1171.32
R73 VSS.n29 VSS 918.774
R74 VSS VSS.t58 918.774
R75 VSS.t48 VSS.t66 826.054
R76 VSS.t41 VSS.t17 826.054
R77 VSS.t25 VSS.t0 792.337
R78 VSS.n150 VSS.n149 767.294
R79 VSS.n169 VSS.n168 767.294
R80 VSS.n157 VSS.n156 763.106
R81 VSS.n177 VSS.n5 763.106
R82 VSS.n150 VSS.n18 732.236
R83 VSS.n168 VSS.n165 732.236
R84 VSS.n157 VSS.n12 732.236
R85 VSS.n181 VSS.n5 732.236
R86 VSS.n29 VSS.n22 708.047
R87 VSS.t46 VSS.t44 708.047
R88 VSS.t62 VSS.t25 708.047
R89 VSS.t5 VSS.t23 708.047
R90 VSS.t51 VSS.t19 708.047
R91 VSS.n93 VSS.t2 681.482
R92 VSS VSS.t46 564.751
R93 VSS VSS.t5 564.751
R94 VSS.t19 VSS 564.751
R95 VSS.n145 VSS 564.751
R96 VSS.t64 VSS.t60 554.492
R97 VSS.t32 VSS.t51 522.606
R98 VSS.t60 VSS.n22 513.419
R99 VSS VSS.t43 480.461
R100 VSS VSS.t20 459.26
R101 VSS.t2 VSS 459.26
R102 VSS.t14 VSS.t64 431.272
R103 VSS.t58 VSS.t32 387.74
R104 VSS.t15 VSS 370.37
R105 VSS.t56 VSS 370.37
R106 VSS.t30 VSS 370.37
R107 VSS VSS.t14 343.991
R108 VSS.n144 VSS.t50 337.166
R109 VSS.n92 VSS.n41 334.815
R110 VSS.n149 VSS.n148 325.502
R111 VSS.n170 VSS.n169 325.502
R112 VSS.t66 VSS.n144 320.307
R113 VSS.n156 VSS.n155 304.204
R114 VSS.n177 VSS.n176 304.204
R115 VSS VSS.t50 295.019
R116 VSS.t20 VSS.n40 278.519
R117 VSS.t0 VSS 261.303
R118 VSS.t10 VSS.t15 248.889
R119 VSS.t54 VSS.t56 248.889
R120 VSS.t35 VSS.t37 248.889
R121 VSS.t28 VSS.t30 248.889
R122 VSS VSS.t7 244.445
R123 VSS.n148 VSS.n21 242.448
R124 VSS.n170 VSS.n162 242.448
R125 VSS.n155 VSS.n15 242.448
R126 VSS.n176 VSS.n4 242.448
R127 VSS.n81 VSS.t1 240.575
R128 VSS.n137 VSS.t13 237.327
R129 VSS.n152 VSS.t27 224.799
R130 VSS.n41 VSS 222.222
R131 VSS.n93 VSS 222.222
R132 VSS.n47 VSS.t68 218.308
R133 VSS.n33 VSS.t71 218.308
R134 VSS.n138 VSS.t69 218.308
R135 VSS.n64 VSS.t70 218.308
R136 VSS.n55 VSS.t3 214.456
R137 VSS.n50 VSS.t4 214.456
R138 VSS.n122 VSS.t21 214.456
R139 VSS.n34 VSS.t22 214.456
R140 VSS.n27 VSS.t8 214.456
R141 VSS.n26 VSS.t9 214.456
R142 VSS.n59 VSS.t33 214.456
R143 VSS.n63 VSS.t34 214.456
R144 VSS.n127 VSS.n126 204.457
R145 VSS.n72 VSS.n71 200.231
R146 VSS.n24 VSS.n23 200.231
R147 VSS.n66 VSS.n61 200.105
R148 VSS VSS.t10 198.519
R149 VSS VSS.t54 198.519
R150 VSS VSS.t35 198.519
R151 VSS VSS.t28 198.519
R152 VSS.n178 VSS.n177 195
R153 VSS.t40 VSS.n178 195
R154 VSS.n180 VSS.n179 195
R155 VSS.n179 VSS.t40 195
R156 VSS.n169 VSS.n161 195
R157 VSS.n161 VSS.t53 195
R158 VSS.n164 VSS.n160 195
R159 VSS.n160 VSS.t53 195
R160 VSS.n156 VSS.n11 195
R161 VSS.n11 VSS.t39 195
R162 VSS.n13 VSS.n10 195
R163 VSS.n10 VSS.t39 195
R164 VSS.n20 VSS.n16 195
R165 VSS.n92 VSS.n16 195
R166 VSS.n149 VSS.n17 195
R167 VSS.n17 VSS.t27 195
R168 VSS.t17 VSS 177.012
R169 VSS.n175 VSS.n6 167.018
R170 VSS.n115 VSS.t16 162.471
R171 VSS.n110 VSS.t57 162.471
R172 VSS.n39 VSS.t38 162.471
R173 VSS.n101 VSS.t31 162.471
R174 VSS.n82 VSS.t26 162.471
R175 VSS.n72 VSS.t24 160.046
R176 VSS.n24 VSS.t45 160.046
R177 VSS.n36 VSS.t11 160.017
R178 VSS.n108 VSS.t55 160.017
R179 VSS.n102 VSS.t36 160.017
R180 VSS.n44 VSS.t29 160.017
R181 VSS.n89 VSS.t6 160.017
R182 VSS.n84 VSS.t63 160.017
R183 VSS.n81 VSS.t47 158.534
R184 VSS.n166 VSS.t53 156.078
R185 VSS.n159 VSS.t39 155.954
R186 VSS.n147 VSS.n146 141.745
R187 VSS VSS.t27 121.481
R188 VSS.n174 VSS.n8 99.9606
R189 VSS.n173 VSS.n172 93.8227
R190 VSS.n153 VSS.n9 93.748
R191 VSS.t37 VSS.n92 85.9264
R192 VSS.t43 VSS.t62 84.2917
R193 VSS.n126 VSS.t65 72.8576
R194 VSS.n61 VSS.t52 72.8576
R195 VSS.n173 VSS.t53 62.2564
R196 VSS.t39 VSS.n9 62.2068
R197 VSS.n71 VSS.t18 58.5719
R198 VSS.n23 VSS.t67 58.5719
R199 VSS.n175 VSS.n174 56.0836
R200 VSS.t44 VSS.t48 50.5752
R201 VSS.t23 VSS.t41 50.5752
R202 VSS.n125 VSS 43.9579
R203 VSS.n128 VSS.n125 34.6358
R204 VSS.n132 VSS.n30 34.6358
R205 VSS.n20 VSS.n18 30.8711
R206 VSS.n165 VSS.n164 30.8711
R207 VSS.n13 VSS.n12 30.8711
R208 VSS.n181 VSS.n180 30.8711
R209 VSS.n94 VSS.n45 26.9246
R210 VSS.n133 VSS.n132 25.6926
R211 VSS.n71 VSS.t42 25.4291
R212 VSS.n23 VSS.t49 25.4291
R213 VSS.n115 VSS.n114 25.224
R214 VSS.n114 VSS.n36 25.224
R215 VSS.n110 VSS.n109 25.224
R216 VSS.n109 VSS.n108 25.224
R217 VSS.n103 VSS.n39 25.224
R218 VSS.n103 VSS.n102 25.224
R219 VSS.n101 VSS.n100 25.224
R220 VSS.n100 VSS.n44 25.224
R221 VSS.n89 VSS.n88 25.224
R222 VSS.n83 VSS.n82 25.224
R223 VSS.n84 VSS.n83 25.224
R224 VSS.n81 VSS.n80 24.0946
R225 VSS.n146 VSS.t27 24.0161
R226 VSS.n126 VSS.t61 22.3257
R227 VSS.n61 VSS.t59 22.3257
R228 VSS.n88 VSS.n72 21.4593
R229 VSS.n80 VSS.n24 21.4593
R230 VSS.n110 VSS.n36 20.3299
R231 VSS.n102 VSS.n101 20.3299
R232 VSS.n116 VSS.n115 19.2926
R233 VSS.n89 VSS.n70 17.7867
R234 VSS.n107 VSS.n39 17.3181
R235 VSS.t7 VSS.t12 16.8587
R236 VSS.n108 VSS.n107 15.8123
R237 VSS.n45 VSS.n44 15.8123
R238 VSS.n56 VSS.n45 14.775
R239 VSS.n143 VSS.n142 14.775
R240 VSS.n82 VSS.n81 13.5534
R241 VSS.n124 VSS.n123 11.2844
R242 VSS.n176 VSS.n7 11.0382
R243 VSS.n8 VSS.n7 11.0382
R244 VSS.n6 VSS.n5 11.0382
R245 VSS.n171 VSS.n170 11.0382
R246 VSS.n172 VSS.n171 11.0382
R247 VSS.n168 VSS.n167 11.0382
R248 VSS.n167 VSS.n166 11.0382
R249 VSS.n155 VSS.n154 11.0382
R250 VSS.n154 VSS.n153 11.0382
R251 VSS.n158 VSS.n157 11.0382
R252 VSS.n159 VSS.n158 11.0382
R253 VSS.n148 VSS.n147 11.0382
R254 VSS.n151 VSS.n150 11.0382
R255 VSS.n152 VSS.n151 11.0382
R256 VSS.n21 VSS.n20 10.9181
R257 VSS.n164 VSS.n162 10.9181
R258 VSS.n15 VSS.n13 10.9181
R259 VSS.n180 VSS.n4 10.9181
R260 VSS.n19 VSS.n18 10.4476
R261 VSS.n165 VSS.n163 10.4476
R262 VSS.n14 VSS.n12 10.4476
R263 VSS.n182 VSS.n181 10.4476
R264 VSS.n84 VSS.n72 10.1652
R265 VSS.n51 VSS.n50 9.70901
R266 VSS.n123 VSS.n122 9.70901
R267 VSS.n63 VSS.n62 9.70901
R268 VSS.n127 VSS.n30 9.41227
R269 VSS.n134 VSS.n133 9.3005
R270 VSS.n136 VSS.n135 9.3005
R271 VSS.n76 VSS.n24 9.3005
R272 VSS.n81 VSS.n75 9.3005
R273 VSS.n86 VSS.n72 9.3005
R274 VSS.n65 VSS.n60 9.3005
R275 VSS.n68 VSS.n67 9.3005
R276 VSS.n70 VSS.n69 9.3005
R277 VSS.n90 VSS.n89 9.3005
R278 VSS.n88 VSS.n87 9.3005
R279 VSS.n85 VSS.n84 9.3005
R280 VSS.n83 VSS.n73 9.3005
R281 VSS.n82 VSS.n74 9.3005
R282 VSS.n80 VSS.n79 9.3005
R283 VSS.n143 VSS.n25 9.3005
R284 VSS.n142 VSS.n141 9.3005
R285 VSS.n140 VSS.n139 9.3005
R286 VSS.n132 VSS.n131 9.3005
R287 VSS.n130 VSS.n30 9.3005
R288 VSS.n129 VSS.n128 9.3005
R289 VSS.n125 VSS.n31 9.3005
R290 VSS.n95 VSS.n94 9.3005
R291 VSS.n98 VSS.n44 9.3005
R292 VSS.n102 VSS.n42 9.3005
R293 VSS.n107 VSS.n106 9.3005
R294 VSS.n108 VSS.n38 9.3005
R295 VSS.n112 VSS.n36 9.3005
R296 VSS.n117 VSS.n116 9.3005
R297 VSS.n120 VSS.n119 9.3005
R298 VSS.n121 VSS.n32 9.3005
R299 VSS.n115 VSS.n35 9.3005
R300 VSS.n114 VSS.n113 9.3005
R301 VSS.n111 VSS.n110 9.3005
R302 VSS.n109 VSS.n37 9.3005
R303 VSS.n105 VSS.n39 9.3005
R304 VSS.n104 VSS.n103 9.3005
R305 VSS.n101 VSS.n43 9.3005
R306 VSS.n100 VSS.n99 9.3005
R307 VSS.n53 VSS.n52 9.3005
R308 VSS.n54 VSS.n46 9.3005
R309 VSS.n57 VSS.n56 9.3005
R310 VSS.n97 VSS.n45 9.3005
R311 VSS.n184 VSS.n183 8.45078
R312 VSS.n186 VSS.n1 8.30267
R313 VSS.n185 VSS.n2 7.97888
R314 VSS.n184 VSS.n3 7.97601
R315 VSS.n19 VSS.n1 7.16724
R316 VSS.n163 VSS.n3 7.16724
R317 VSS.n14 VSS.n2 7.16724
R318 VSS.n183 VSS.n182 7.16724
R319 VSS.n143 VSS.n24 7.15344
R320 VSS.n96 VSS.n91 6.50373
R321 VSS.n128 VSS.n127 6.4005
R322 VSS.n54 VSS.n53 6.26433
R323 VSS.n121 VSS.n120 6.26433
R324 VSS.n55 VSS.n54 5.85582
R325 VSS.n122 VSS.n121 5.85582
R326 VSS.n67 VSS.n59 5.85582
R327 VSS.n136 VSS.n27 5.85582
R328 VSS.n139 VSS.n137 5.85582
R329 VSS.n97 VSS.n96 4.788
R330 VSS.n21 VSS.n19 4.73093
R331 VSS.n163 VSS.n162 4.73093
R332 VSS.n15 VSS.n14 4.73093
R333 VSS.n182 VSS.n4 4.73093
R334 VSS.n96 VSS.n95 4.50726
R335 VSS.n187 VSS 4.01425
R336 VSS.n66 VSS.n65 3.40476
R337 VSS.n53 VSS.n47 3.13241
R338 VSS.n120 VSS.n33 3.13241
R339 VSS.n65 VSS.n64 3.13241
R340 VSS.n139 VSS.n138 3.13241
R341 VSS.n77 VSS.n28 2.88636
R342 VSS.n67 VSS.n66 2.86007
R343 VSS.n50 VSS.n47 2.7239
R344 VSS.n34 VSS.n33 2.7239
R345 VSS.n64 VSS.n63 2.7239
R346 VSS.n138 VSS.n26 2.7239
R347 VSS.n118 VSS.n0 1.753
R348 VSS.n49 VSS.n48 1.753
R349 VSS.n78 VSS.n77 1.21169
R350 VSS.n48 VSS.n0 0.761313
R351 VSS.n188 VSS.n0 0.591917
R352 VSS.n77 VSS 0.531208
R353 VSS.n188 VSS.n187 0.506165
R354 VSS.n185 VSS.n184 0.467019
R355 VSS.n56 VSS.n55 0.409011
R356 VSS.n116 VSS.n34 0.409011
R357 VSS.n70 VSS.n59 0.409011
R358 VSS.n133 VSS.n27 0.409011
R359 VSS.n137 VSS.n136 0.409011
R360 VSS.n142 VSS.n26 0.409011
R361 VSS.n187 VSS.n186 0.198729
R362 VSS.n95 VSS.n58 0.1255
R363 VSS.n129 VSS.n31 0.120292
R364 VSS.n130 VSS.n129 0.120292
R365 VSS.n131 VSS.n130 0.120292
R366 VSS.n141 VSS.n140 0.120292
R367 VSS.n74 VSS.n73 0.120292
R368 VSS.n85 VSS.n73 0.120292
R369 VSS.n87 VSS.n86 0.120292
R370 VSS.n69 VSS.n68 0.120292
R371 VSS.n68 VSS.n60 0.120292
R372 VSS.n62 VSS.n60 0.120292
R373 VSS.n123 VSS.n32 0.120292
R374 VSS.n119 VSS.n32 0.120292
R375 VSS.n113 VSS.n35 0.120292
R376 VSS.n113 VSS.n112 0.120292
R377 VSS.n111 VSS.n37 0.120292
R378 VSS.n38 VSS.n37 0.120292
R379 VSS.n105 VSS.n104 0.120292
R380 VSS.n104 VSS.n42 0.120292
R381 VSS.n99 VSS.n43 0.120292
R382 VSS.n99 VSS.n98 0.120292
R383 VSS.n57 VSS.n46 0.120292
R384 VSS.n52 VSS.n51 0.120292
R385 VSS.n140 VSS 0.0981562
R386 VSS VSS.n124 0.09425
R387 VSS.n48 VSS 0.0881354
R388 VSS.n186 VSS.n185 0.0766574
R389 VSS.n52 VSS.n49 0.0721146
R390 VSS.n79 VSS.n78 0.0708125
R391 VSS.n1 VSS 0.064875
R392 VSS.n3 VSS 0.064875
R393 VSS.n2 VSS 0.064875
R394 VSS.n183 VSS 0.063625
R395 VSS.n119 VSS.n118 0.0616979
R396 VSS.n131 VSS 0.0603958
R397 VSS.n135 VSS 0.0603958
R398 VSS VSS.n25 0.0603958
R399 VSS.n76 VSS 0.0603958
R400 VSS.n79 VSS 0.0603958
R401 VSS VSS.n75 0.0603958
R402 VSS VSS.n74 0.0603958
R403 VSS.n86 VSS 0.0603958
R404 VSS.n87 VSS 0.0603958
R405 VSS.n69 VSS 0.0603958
R406 VSS.n35 VSS 0.0603958
R407 VSS VSS.n111 0.0603958
R408 VSS.n106 VSS 0.0603958
R409 VSS VSS.n105 0.0603958
R410 VSS.n43 VSS 0.0603958
R411 VSS VSS.n97 0.0603958
R412 VSS VSS.n57 0.0603958
R413 VSS.n91 VSS 0.0590938
R414 VSS.n118 VSS.n117 0.0590938
R415 VSS.n78 VSS.n76 0.0499792
R416 VSS.n49 VSS.n46 0.0486771
R417 VSS VSS.n28 0.0460729
R418 VSS VSS.n134 0.0343542
R419 VSS VSS.n25 0.0330521
R420 VSS.n106 VSS 0.0330521
R421 VSS.n58 VSS 0.03175
R422 VSS VSS.n188 0.0292529
R423 VSS.t40 VSS.n175 0.0270008
R424 VSS.n135 VSS 0.0226354
R425 VSS.n141 VSS 0.0226354
R426 VSS.n75 VSS 0.0226354
R427 VSS VSS.n85 0.0226354
R428 VSS.n90 VSS 0.0226354
R429 VSS.n62 VSS 0.0226354
R430 VSS.n117 VSS 0.0226354
R431 VSS.n112 VSS 0.0226354
R432 VSS VSS.n38 0.0226354
R433 VSS VSS.n42 0.0226354
R434 VSS.n98 VSS 0.0226354
R435 VSS.n51 VSS 0.0226354
R436 VSS.n134 VSS.n28 0.0148229
R437 VSS.n124 VSS.n31 0.00440625
R438 VSS.n91 VSS.n90 0.00180208
R439 VSS.n97 VSS.n58 0.00180208
R440 VDD.n177 VDD.n175 8629.41
R441 VDD.n180 VDD.n174 8629.41
R442 VDD.n161 VDD.n160 8629.41
R443 VDD.n163 VDD.n158 8629.41
R444 VDD.n144 VDD.n143 8629.41
R445 VDD.n146 VDD.n141 8629.41
R446 VDD.n127 VDD.n125 8629.41
R447 VDD.n130 VDD.n124 8629.41
R448 VDD.n176 VDD.n173 920.471
R449 VDD.n164 VDD.n157 920.471
R450 VDD.n147 VDD.n140 920.471
R451 VDD.n126 VDD.n123 920.471
R452 VDD.n182 VDD.n173 914.447
R453 VDD.n166 VDD.n164 914.447
R454 VDD.n149 VDD.n147 914.447
R455 VDD.n132 VDD.n123 914.447
R456 VDD.t7 VDD.n59 804.731
R457 VDD.n61 VDD.t7 751.692
R458 VDD.n33 VDD.t64 671.408
R459 VDD.n22 VDD.t27 671.408
R460 VDD VDD.t6 630.375
R461 VDD.n92 VDD.n91 602.456
R462 VDD.n114 VDD.n2 602.456
R463 VDD.n6 VDD.n5 585
R464 VDD.n8 VDD.n7 585
R465 VDD.n176 VDD.n120 480.764
R466 VDD.n157 VDD.n155 480.764
R467 VDD.n140 VDD.n138 480.764
R468 VDD.n126 VDD.n122 480.764
R469 VDD VDD.t9 458.724
R470 VDD.t6 VDD 458.724
R471 VDD.n54 VDD.t41 420.25
R472 VDD.n50 VDD.t10 388.656
R473 VDD.n85 VDD.t11 388.656
R474 VDD.n63 VDD.t8 388.656
R475 VDD.n36 VDD.t4 388.656
R476 VDD.n45 VDD.t5 388.656
R477 VDD.n10 VDD.t13 388.656
R478 VDD.n15 VDD.t14 388.656
R479 VDD.n184 VDD.n120 379.2
R480 VDD.n168 VDD.n155 379.2
R481 VDD.n151 VDD.n138 379.2
R482 VDD.n134 VDD.n122 379.2
R483 VDD VDD.t15 369.938
R484 VDD VDD.t67 369.938
R485 VDD.n39 VDD.n32 322.329
R486 VDD.n17 VDD.n13 322.329
R487 VDD.n96 VDD.n94 259.697
R488 VDD.n72 VDD.t68 255.905
R489 VDD.n77 VDD.t16 255.905
R490 VDD.n53 VDD.t42 255.905
R491 VDD.n93 VDD.t52 255.905
R492 VDD.n43 VDD.t23 254.475
R493 VDD.n68 VDD.t18 252.95
R494 VDD.n73 VDD.t70 252.95
R495 VDD.n78 VDD.t44 252.95
R496 VDD.n113 VDD.t34 252.95
R497 VDD.n92 VDD.t60 251.516
R498 VDD.n3 VDD.t32 250.724
R499 VDD.n1 VDD.t36 250.724
R500 VDD.t41 VDD.t43 248.599
R501 VDD.t15 VDD.t69 248.599
R502 VDD.t67 VDD.t17 248.599
R503 VDD.n108 VDD.t30 248.219
R504 VDD.n95 VDD.t54 248.219
R505 VDD.n54 VDD 221.964
R506 VDD.n61 VDD.t74 215.827
R507 VDD.n43 VDD.n42 213.119
R508 VDD.n83 VDD.n54 213.119
R509 VDD.n51 VDD.t72 210.964
R510 VDD.n37 VDD.t73 210.964
R511 VDD.n12 VDD.t71 210.964
R512 VDD.n103 VDD.n102 209.368
R513 VDD.t43 VDD 198.287
R514 VDD.t69 VDD 198.287
R515 VDD.t17 VDD 198.287
R516 VDD.n105 VDD.n104 183.673
R517 VDD VDD.t61 182.952
R518 VDD VDD.n103 182.952
R519 VDD.t55 VDD 182.952
R520 VDD.n7 VDD.n6 159.476
R521 VDD.n94 VDD.t2 157.014
R522 VDD.t31 VDD.t19 154.417
R523 VDD.t47 VDD.t1 147.703
R524 VDD.t65 VDD.t63 140.989
R525 VDD.t1 VDD.t53 140.989
R526 VDD.t33 VDD.t35 140.989
R527 VDD.t29 VDD.t31 140.989
R528 VDD.t26 VDD.t49 140.989
R529 VDD.n94 VDD.t46 137.079
R530 VDD.n42 VDD 125.883
R531 VDD.n104 VDD 125.883
R532 VDD.n32 VDD.t66 116.341
R533 VDD.n13 VDD.t50 116.341
R534 VDD.t63 VDD 112.457
R535 VDD.t53 VDD 112.457
R536 VDD VDD.t26 112.457
R537 VDD VDD.t37 109.1
R538 VDD.t3 VDD.t65 104.064
R539 VDD.t49 VDD.t12 104.064
R540 VDD.t24 VDD 102.385
R541 VDD.t22 VDD 99.0288
R542 VDD.n91 VDD.t48 96.1553
R543 VDD.n2 VDD.t40 96.1553
R544 VDD VDD.t39 92.315
R545 VDD.n6 VDD.t20 86.7743
R546 VDD.n42 VDD.t22 83.9228
R547 VDD.n103 VDD.t45 80.5659
R548 VDD.t61 VDD.t3 77.209
R549 VDD.t12 VDD.t55 77.209
R550 VDD.n7 VDD.t38 66.8398
R551 VDD.n183 VDD.n182 66.6358
R552 VDD.n167 VDD.n166 66.6358
R553 VDD.n150 VDD.n149 66.6358
R554 VDD.n133 VDD.n132 66.6358
R555 VDD.n91 VDD.t25 63.3219
R556 VDD.n2 VDD.t58 63.3219
R557 VDD VDD.t47 62.103
R558 VDD.n177 VDD.n176 61.6672
R559 VDD.n181 VDD.n180 61.6672
R560 VDD.n161 VDD.n157 61.6672
R561 VDD.n158 VDD.n156 61.6672
R562 VDD.n144 VDD.n140 61.6672
R563 VDD.n141 VDD.n139 61.6672
R564 VDD.n127 VDD.n126 61.6672
R565 VDD.n131 VDD.n130 61.6672
R566 VDD.n178 VDD.n177 60.9564
R567 VDD.n180 VDD.n179 60.9564
R568 VDD.n162 VDD.n161 60.9564
R569 VDD.n159 VDD.n158 60.9564
R570 VDD.n145 VDD.n144 60.9564
R571 VDD.n142 VDD.n141 60.9564
R572 VDD.n128 VDD.n127 60.9564
R573 VDD.n130 VDD.n129 60.9564
R574 VDD.n167 VDD.n156 60.6123
R575 VDD.n150 VDD.n139 60.6123
R576 VDD.n183 VDD.n172 59.4829
R577 VDD.n133 VDD.n121 58.7299
R578 VDD.t19 VDD 55.3892
R579 VDD.t57 VDD 52.0323
R580 VDD VDD.t45 45.3185
R581 VDD VDD.t59 41.9616
R582 VDD.n178 VDD.n174 38.5759
R583 VDD.n179 VDD.n175 38.5759
R584 VDD.n163 VDD.n162 38.5759
R585 VDD.n160 VDD.n159 38.5759
R586 VDD.n146 VDD.n145 38.5759
R587 VDD.n143 VDD.n142 38.5759
R588 VDD.n128 VDD.n124 38.5759
R589 VDD.n129 VDD.n125 38.5759
R590 VDD.n102 VDD.n24 34.6358
R591 VDD.n102 VDD.n25 34.6358
R592 VDD.n107 VDD.n106 34.6358
R593 VDD.n104 VDD 28.5341
R594 VDD.n32 VDD.t62 28.4453
R595 VDD.n13 VDD.t56 28.4453
R596 VDD.n109 VDD.n108 28.3534
R597 VDD.n106 VDD.n105 25.6953
R598 VDD.n72 VDD.n57 25.224
R599 VDD.n68 VDD.n57 25.224
R600 VDD.n77 VDD.n56 25.224
R601 VDD.n73 VDD.n56 25.224
R602 VDD.n79 VDD.n53 25.224
R603 VDD.n79 VDD.n78 25.224
R604 VDD.n97 VDD.n93 25.224
R605 VDD.n43 VDD.n27 23.7181
R606 VDD VDD.n33 23.252
R607 VDD.n92 VDD.n27 21.4593
R608 VDD.n73 VDD.n72 20.3299
R609 VDD.n78 VDD.n77 20.3299
R610 VDD.t39 VDD.t33 20.1418
R611 VDD.n114 VDD.n1 19.9534
R612 VDD.n113 VDD.n112 19.8181
R613 VDD.n83 VDD.n53 17.3181
R614 VDD.n96 VDD.n95 17.3181
R615 VDD.n93 VDD.n92 16.5652
R616 VDD.n97 VDD.n96 16.5652
R617 VDD.n68 VDD.n67 15.8123
R618 VDD.n84 VDD.n83 14.2735
R619 VDD.n44 VDD.n43 14.2735
R620 VDD.n106 VDD.n22 13.9299
R621 VDD.n119 VDD.n118 13.6791
R622 VDD.n114 VDD.n113 13.5534
R623 VDD.n49 VDD.n48 11.4366
R624 VDD.n185 VDD.n184 11.3235
R625 VDD.n169 VDD.n168 11.3235
R626 VDD.n152 VDD.n151 11.3235
R627 VDD.n135 VDD.n134 11.3235
R628 VDD.n105 VDD.n23 11.2937
R629 VDD.n89 VDD.n88 11.2737
R630 VDD.t59 VDD.t24 10.0712
R631 VDD.n63 VDD.n60 9.60526
R632 VDD.n50 VDD.n49 9.60526
R633 VDD.n15 VDD.n14 9.60526
R634 VDD.n52 VDD.n28 9.3005
R635 VDD.n87 VDD.n86 9.3005
R636 VDD.n84 VDD.n29 9.3005
R637 VDD.n83 VDD.n82 9.3005
R638 VDD.n78 VDD.n55 9.3005
R639 VDD.n74 VDD.n73 9.3005
R640 VDD.n69 VDD.n68 9.3005
R641 VDD.n65 VDD.n64 9.3005
R642 VDD.n70 VDD.n57 9.3005
R643 VDD.n72 VDD.n71 9.3005
R644 VDD.n75 VDD.n56 9.3005
R645 VDD.n77 VDD.n76 9.3005
R646 VDD.n80 VDD.n79 9.3005
R647 VDD.n81 VDD.n53 9.3005
R648 VDD.n110 VDD.n109 9.3005
R649 VDD.n115 VDD.n114 9.3005
R650 VDD.n99 VDD.n24 9.3005
R651 VDD.n92 VDD.n90 9.3005
R652 VDD.n43 VDD.n41 9.3005
R653 VDD.n35 VDD.n34 9.3005
R654 VDD.n38 VDD.n30 9.3005
R655 VDD.n47 VDD.n46 9.3005
R656 VDD.n44 VDD.n31 9.3005
R657 VDD.n40 VDD.n27 9.3005
R658 VDD.n93 VDD.n26 9.3005
R659 VDD.n98 VDD.n97 9.3005
R660 VDD.n102 VDD.n101 9.3005
R661 VDD.n100 VDD.n25 9.3005
R662 VDD.n113 VDD.n0 9.3005
R663 VDD.n112 VDD.n111 9.3005
R664 VDD.n107 VDD.n4 9.3005
R665 VDD.n106 VDD.n9 9.3005
R666 VDD.n21 VDD.n20 9.3005
R667 VDD.n19 VDD.n18 9.3005
R668 VDD.n16 VDD.n11 9.3005
R669 VDD.n136 VDD.n121 8.23557
R670 VDD.n8 VDD.n5 6.8005
R671 VDD.n67 VDD.n59 6.48583
R672 VDD.n182 VDD.n181 6.02403
R673 VDD.n132 VDD.n131 6.02403
R674 VDD.n62 VDD.n61 5.8885
R675 VDD.n165 VDD.n156 4.89462
R676 VDD.n149 VDD.n148 4.89462
R677 VDD.n86 VDD.n52 4.67352
R678 VDD.n67 VDD.n66 4.62124
R679 VDD.n64 VDD.n63 4.36875
R680 VDD.n86 VDD.n85 4.36875
R681 VDD.n46 VDD.n45 4.36875
R682 VDD.n16 VDD.n15 4.36875
R683 VDD.t35 VDD.t57 3.35739
R684 VDD.t37 VDD.t29 3.35739
R685 VDD.n165 VDD.n154 3.23917
R686 VDD.n148 VDD.n137 3.23136
R687 VDD.n172 VDD.n171 3.22655
R688 VDD.n64 VDD.n62 3.2005
R689 VDD.n174 VDD.n173 2.84665
R690 VDD.n175 VDD.n120 2.84665
R691 VDD.n164 VDD.n163 2.84665
R692 VDD.n160 VDD.n155 2.84665
R693 VDD.n147 VDD.n146 2.84665
R694 VDD.n143 VDD.n138 2.84665
R695 VDD.n124 VDD.n123 2.84665
R696 VDD.n125 VDD.n122 2.84665
R697 VDD.n62 VDD.n59 2.8165
R698 VDD.n39 VDD.n38 2.54018
R699 VDD.n18 VDD.n17 2.54018
R700 VDD.n52 VDD.n51 2.33701
R701 VDD.n38 VDD.n37 2.33701
R702 VDD.n18 VDD.n12 2.33701
R703 VDD.n184 VDD.n183 2.28169
R704 VDD.n168 VDD.n167 2.28169
R705 VDD.n151 VDD.n150 2.28169
R706 VDD.n134 VDD.n133 2.28169
R707 VDD.n46 VDD.n39 2.13383
R708 VDD.n17 VDD.n16 2.13383
R709 VDD.n51 VDD.n50 2.03225
R710 VDD.n37 VDD.n36 2.03225
R711 VDD.n12 VDD.n10 2.03225
R712 VDD.n131 VDD.n121 1.88285
R713 VDD.n117 VDD.n116 1.753
R714 VDD.n25 VDD.n1 1.50638
R715 VDD.n109 VDD.n8 1.4005
R716 VDD.n35 VDD.n33 1.37193
R717 VDD.n22 VDD.n21 1.37193
R718 VDD.n170 VDD.n169 1.143
R719 VDD.n153 VDD.n152 1.143
R720 VDD.n185 VDD.n119 1.13925
R721 VDD.n136 VDD.n135 1.13675
R722 VDD.n181 VDD.n172 1.12991
R723 VDD.n166 VDD.n165 1.12991
R724 VDD.n148 VDD.n139 1.12991
R725 VDD.n58 VDD 1.06099
R726 VDD.n154 VDD.n153 0.862816
R727 VDD.n137 VDD.n136 0.770881
R728 VDD.n95 VDD.n24 0.753441
R729 VDD.n108 VDD.n107 0.753441
R730 VDD.n171 VDD.n170 0.729231
R731 VDD.n5 VDD.n3 0.6005
R732 VDD.n118 VDD.n117 0.511794
R733 VDD.n117 VDD 0.460219
R734 VDD.n171 VDD.n119 0.405788
R735 VDD.n112 VDD.n3 0.4005
R736 VDD.n153 VDD.n137 0.392323
R737 VDD.n170 VDD.n154 0.360318
R738 VDD.n85 VDD.n84 0.305262
R739 VDD.n36 VDD.n35 0.305262
R740 VDD.n45 VDD.n44 0.305262
R741 VDD.n21 VDD.n10 0.305262
R742 VDD.t28 VDD.n178 0.27666
R743 VDD.n179 VDD.t28 0.27666
R744 VDD.n162 VDD.t0 0.27666
R745 VDD.n159 VDD.t0 0.27666
R746 VDD.n145 VDD.t51 0.27666
R747 VDD.n142 VDD.t51 0.27666
R748 VDD.t21 VDD.n128 0.27666
R749 VDD.n129 VDD.t21 0.27666
R750 VDD.n66 VDD.n65 0.180304
R751 VDD.n66 VDD 0.120408
R752 VDD.n49 VDD.n28 0.120292
R753 VDD.n87 VDD.n29 0.120292
R754 VDD.n81 VDD.n80 0.120292
R755 VDD.n80 VDD.n55 0.120292
R756 VDD.n76 VDD.n75 0.120292
R757 VDD.n75 VDD.n74 0.120292
R758 VDD.n71 VDD.n70 0.120292
R759 VDD.n70 VDD.n69 0.120292
R760 VDD.n65 VDD.n60 0.120292
R761 VDD.n34 VDD.n30 0.120292
R762 VDD.n47 VDD.n31 0.120292
R763 VDD.n98 VDD.n26 0.120292
R764 VDD.n99 VDD.n98 0.120292
R765 VDD.n115 VDD.n0 0.120292
R766 VDD.n111 VDD.n110 0.120292
R767 VDD.n110 VDD.n4 0.120292
R768 VDD.n20 VDD.n19 0.120292
R769 VDD.n19 VDD.n11 0.120292
R770 VDD.n14 VDD.n11 0.120292
R771 VDD.n88 VDD.n28 0.11899
R772 VDD.n34 VDD 0.0981562
R773 VDD.n89 VDD 0.0955521
R774 VDD.n48 VDD.n30 0.0916458
R775 VDD.n169 VDD 0.06425
R776 VDD.n152 VDD 0.06425
R777 VDD.n135 VDD 0.06425
R778 VDD VDD.n185 0.06425
R779 VDD.n82 VDD 0.0603958
R780 VDD VDD.n81 0.0603958
R781 VDD.n76 VDD 0.0603958
R782 VDD.n71 VDD 0.0603958
R783 VDD.n41 VDD 0.0603958
R784 VDD VDD.n40 0.0603958
R785 VDD VDD.n26 0.0603958
R786 VDD.n101 VDD 0.0603958
R787 VDD VDD.n100 0.0603958
R788 VDD.n111 VDD 0.0603958
R789 VDD.n20 VDD 0.0603958
R790 VDD.n23 VDD 0.0590938
R791 VDD.n116 VDD 0.0525833
R792 VDD.n116 VDD.n115 0.0460729
R793 VDD.n41 VDD 0.0382604
R794 VDD VDD.n58 0.0369583
R795 VDD.n82 VDD 0.03175
R796 VDD.n101 VDD 0.03175
R797 VDD.n48 VDD.n47 0.0291458
R798 VDD.n118 VDD 0.0236148
R799 VDD VDD.n29 0.0226354
R800 VDD VDD.n55 0.0226354
R801 VDD.n74 VDD 0.0226354
R802 VDD.n69 VDD 0.0226354
R803 VDD.n60 VDD 0.0226354
R804 VDD VDD.n31 0.0226354
R805 VDD.n40 VDD 0.0226354
R806 VDD.n90 VDD 0.0226354
R807 VDD VDD.n99 0.0226354
R808 VDD.n100 VDD 0.0226354
R809 VDD VDD.n0 0.0226354
R810 VDD VDD.n4 0.0226354
R811 VDD VDD.n9 0.0226354
R812 VDD.n14 VDD 0.0226354
R813 VDD.n90 VDD.n89 0.00310417
R814 VDD.n88 VDD.n87 0.00180208
R815 VDD.n58 VDD 0.00180208
R816 VDD.n23 VDD.n9 0.00180208
R817 A3.n1 A3.t1 26.3998
R818 A3.n1 A3.t0 23.5483
R819 A3.n0 A3.t2 12.7127
R820 A3.n0 A3.t3 10.8578
R821 A3.n2 A3.n1 3.12177
R822 A3.n2 A3.n0 1.81453
R823 A3.n3 A3.n2 1.1255
R824 A3.n3 A3 0.210543
R825 A3 A3.n3 0.0655
R826 Z.n18 Z.t1 23.6581
R827 Z.n12 Z.t11 23.6581
R828 Z.n6 Z.t0 23.6581
R829 Z.n1 Z.t4 23.6581
R830 Z.n20 Z.t2 23.3739
R831 Z.n14 Z.t10 23.3739
R832 Z.n8 Z.t14 23.3739
R833 Z.n3 Z.t3 23.3739
R834 Z.n18 Z.t9 10.7528
R835 Z.n12 Z.t12 10.7528
R836 Z.n6 Z.t7 10.7528
R837 Z.n1 Z.t5 10.7528
R838 Z.n17 Z.t15 10.6417
R839 Z.n11 Z.t13 10.6417
R840 Z.n5 Z.t8 10.6417
R841 Z.n0 Z.t6 10.6417
R842 Z.n19 Z.n18 1.30064
R843 Z.n13 Z.n12 1.30064
R844 Z.n7 Z.n6 1.30064
R845 Z.n2 Z.n1 1.30064
R846 Z Z.n4 0.983856
R847 Z.n22 Z.n21 0.956356
R848 Z.n10 Z.n9 0.936641
R849 Z.n16 Z.n15 0.924585
R850 Z Z.n24 0.753
R851 Z.n20 Z.n19 0.726502
R852 Z.n14 Z.n13 0.726502
R853 Z.n8 Z.n7 0.726502
R854 Z.n3 Z.n2 0.726502
R855 Z.n23 Z 0.723
R856 Z.n19 Z.n17 0.512491
R857 Z.n13 Z.n11 0.512491
R858 Z.n7 Z.n5 0.512491
R859 Z.n2 Z.n0 0.512491
R860 Z Z.n23 0.4155
R861 Z.n21 Z.n17 0.359663
R862 Z.n15 Z.n11 0.359663
R863 Z.n9 Z.n5 0.359663
R864 Z.n4 Z.n0 0.359663
R865 Z.n24 Z 0.25425
R866 Z.n21 Z.n20 0.216071
R867 Z.n15 Z.n14 0.216071
R868 Z.n9 Z.n8 0.216071
R869 Z.n4 Z.n3 0.216071
R870 Z.n24 Z 0.088
R871 Z.n10 Z 0.0776605
R872 Z.n16 Z 0.0656042
R873 Z.n23 Z 0.0655
R874 Z Z.n10 0.0561931
R875 Z Z.n16 0.0376287
R876 Z.n22 Z 0.028
R877 Z Z.n22 0.0274608
R878 mux4onehot_0.x2.GP2.n4 mux4onehot_0.x2.GP2.t4 450.938
R879 mux4onehot_0.x2.GP2.n4 mux4onehot_0.x2.GP2.t5 445.666
R880 mux4onehot_0.x2.GP2.n5 mux4onehot_0.x2.GP2.n3 195.958
R881 mux4onehot_0.x2.GP2.n1 mux4onehot_0.x2.GP2.n0 101.49
R882 mux4onehot_0.x2.GP2.n3 mux4onehot_0.x2.GP2.t3 26.5955
R883 mux4onehot_0.x2.GP2.n3 mux4onehot_0.x2.GP2.t2 26.5955
R884 mux4onehot_0.x2.GP2.n0 mux4onehot_0.x2.GP2.t1 24.9236
R885 mux4onehot_0.x2.GP2.n0 mux4onehot_0.x2.GP2.t0 24.9236
R886 mux4onehot_0.x1.gpo1 mux4onehot_0.x2.x2.GP 13.129
R887 mux4onehot_0.x2.GP2.n5 mux4onehot_0.x1.gpo1 11.995
R888 mux4onehot_0.x2.GP2.n2 mux4onehot_0.x1.x12.Y 10.7525
R889 mux4onehot_0.x1.x12.Y mux4onehot_0.x2.GP2.n5 7.96524
R890 mux4onehot_0.x2.GP2.n2 mux4onehot_0.x1.x12.Y 6.6565
R891 mux4onehot_0.x1.x12.Y mux4onehot_0.x2.GP2.n2 5.04292
R892 mux4onehot_0.x2.x2.GP mux4onehot_0.x2.GP2.n4 2.94361
R893 mux4onehot_0.x1.x12.Y mux4onehot_0.x2.GP2.n1 2.5605
R894 mux4onehot_0.x2.GP2.n1 mux4onehot_0.x1.x12.Y 1.93989
R895 select1.n10 select1.t8 327.99
R896 select1.n3 select1.t0 293.969
R897 select1.n6 select1.t5 256.07
R898 select1.n1 select1.t6 212.081
R899 select1.n0 select1.t3 212.081
R900 select1.n10 select1.t1 199.457
R901 select1.n2 select1.n1 182.929
R902 select1 select1.n3 154.065
R903 select1.n11 select1.n10 152
R904 select1.n7 select1.n6 152
R905 select1.n6 select1.t7 150.03
R906 select1.n1 select1.t4 139.78
R907 select1.n0 select1.t2 139.78
R908 select1.n3 select1.t9 138.338
R909 select1.n1 select1.n0 61.346
R910 select1.n5 select1 22.1096
R911 select1.n14 select1.n13 14.6836
R912 select1.n13 select1.n12 14.6704
R913 select1.n12 select1 13.8672
R914 select1.n4 select1 13.8328
R915 select1.n11 select1 12.1605
R916 select1.n14 select1.n2 10.6811
R917 select1.n7 select1.n5 10.4374
R918 select1.n9 select1.n8 8.15359
R919 select1.n2 select1 6.1445
R920 select1.n4 select1 5.16179
R921 select1.n9 select1.n4 4.65206
R922 select1.n8 select1 3.93896
R923 select1 select1.n11 2.34717
R924 select1.n5 select1 2.16665
R925 select1.n8 select1.n7 1.57588
R926 select1.n13 select1.n9 0.79438
R927 select1.n12 select1 0.6405
R928 select1 select1.n14 0.248606
R929 mux4onehot_0.x2.GP4.n2 mux4onehot_0.x2.GP4.t5 450.938
R930 mux4onehot_0.x2.GP4.n2 mux4onehot_0.x2.GP4.t4 445.666
R931 mux4onehot_0.x1.x14.Y mux4onehot_0.x2.GP4.n4 203.923
R932 mux4onehot_0.x2.GP4.n0 mux4onehot_0.x2.GP4.n1 101.49
R933 mux4onehot_0.x2.GP4.n4 mux4onehot_0.x2.GP4.t2 26.5955
R934 mux4onehot_0.x2.GP4.n4 mux4onehot_0.x2.GP4.t3 26.5955
R935 mux4onehot_0.x2.GP4.n1 mux4onehot_0.x2.GP4.t1 24.9236
R936 mux4onehot_0.x2.GP4.n1 mux4onehot_0.x2.GP4.t0 24.9236
R937 mux4onehot_0.x1.gpo3 mux4onehot_0.x2.x4.GP 16.5752
R938 mux4onehot_0.x2.GP4.n3 mux4onehot_0.x1.x14.Y 10.7525
R939 mux4onehot_0.x2.GP4.n0 mux4onehot_0.x1.gpo3 7.7042
R940 mux4onehot_0.x2.GP4.n3 mux4onehot_0.x1.x14.Y 6.6565
R941 mux4onehot_0.x1.x14.Y mux4onehot_0.x2.GP4.n3 5.04292
R942 mux4onehot_0.x2.x4.GP mux4onehot_0.x2.GP4.n2 2.95993
R943 mux4onehot_0.x1.x14.Y mux4onehot_0.x2.GP4.n0 2.5605
R944 mux4onehot_0.x2.GP4.n0 mux4onehot_0.x1.x14.Y 1.93989
R945 A4.n1 A4.t1 26.3998
R946 A4.n1 A4.t2 23.5483
R947 A4.n0 A4.t3 12.7127
R948 A4.n0 A4.t0 10.8578
R949 A4.n2 A4.n1 3.12177
R950 A4.n2 A4.n0 1.81453
R951 A4.n3 A4.n2 1.1255
R952 A4 A4.n3 0.203263
R953 A4.n3 A4 0.0655
R954 mux4onehot_0.x2.GN4.n1 mux4onehot_0.x2.GN4.t6 377.486
R955 mux4onehot_0.x2.GN4.n1 mux4onehot_0.x2.GN4.t4 374.202
R956 mux4onehot_0.x2.GN4.n7 mux4onehot_0.x2.GN4.t1 339.418
R957 mux4onehot_0.x2.GN4.n0 mux4onehot_0.x2.GN4.t0 274.06
R958 mux4onehot_0.x2.GN4.n4 mux4onehot_0.x2.GN4.t3 212.081
R959 mux4onehot_0.x2.GN4.n3 mux4onehot_0.x2.GN4.t2 212.081
R960 mux4onehot_0.x2.GN4.n5 mux4onehot_0.x2.GN4.n4 184.977
R961 mux4onehot_0.x2.GN4.n4 mux4onehot_0.x2.GN4.t7 139.78
R962 mux4onehot_0.x2.GN4.n3 mux4onehot_0.x2.GN4.t5 139.78
R963 mux4onehot_0.x2.GN4.n4 mux4onehot_0.x2.GN4.n3 61.346
R964 mux4onehot_0.x2.GN4.n6 mux4onehot_0.x2.GN4 18.2601
R965 mux4onehot_0.x2.GN4 mux4onehot_0.x2.GN4.n2 17.2682
R966 mux4onehot_0.x2.GN4 mux4onehot_0.x2.GN4.n5 15.0136
R967 mux4onehot_0.x2.GN4 mux4onehot_0.x2.GN4.n0 11.2645
R968 mux4onehot_0.x2.GN4 mux4onehot_0.x2.GN4.n6 8.9605
R969 mux4onehot_0.x2.GN4.n6 mux4onehot_0.x2.GN4 8.4485
R970 mux4onehot_0.x2.GN4.n2 mux4onehot_0.x2.GN4 8.19806
R971 mux4onehot_0.x2.GN4.n8 mux4onehot_0.x2.GN4 6.6565
R972 mux4onehot_0.x2.GN4.n0 mux4onehot_0.x2.GN4 6.1445
R973 mux4onehot_0.x2.GN4.n2 mux4onehot_0.x2.GN4 4.58237
R974 mux4onehot_0.x2.GN4.n5 mux4onehot_0.x2.GN4 4.0965
R975 mux4onehot_0.x2.GN4.n8 mux4onehot_0.x2.GN4.n7 4.0914
R976 mux4onehot_0.x2.GN4 mux4onehot_0.x2.GN4.n8 3.61789
R977 mux4onehot_0.x2.GN4.n0 mux4onehot_0.x2.GN4 2.86947
R978 mux4onehot_0.x2.GN4 mux4onehot_0.x2.GN4.n1 2.04102
R979 mux4onehot_0.x2.GN4.n7 mux4onehot_0.x2.GN4 1.74382
R980 nselect2.n5 nselect2.n4 196.339
R981 nselect2.n1 nselect2.n0 101.49
R982 nselect2.n4 nselect2.t2 26.5955
R983 nselect2.n4 nselect2.t3 26.5955
R984 nselect2.n0 nselect2.t0 24.9236
R985 nselect2.n0 nselect2.t1 24.9236
R986 nselect2.n2 nselect2 13.5685
R987 nselect2.n3 nselect2 10.7525
R988 nselect2.n6 nselect2.n2 9.50196
R989 nselect2.n6 nselect2.n5 7.64514
R990 nselect2.n5 nselect2 7.58449
R991 nselect2.n3 nselect2 6.6565
R992 nselect2 nselect2.n3 5.04292
R993 nselect2 nselect2.n2 3.8405
R994 nselect2 nselect2.n1 2.5605
R995 nselect2.n1 nselect2 1.93989
R996 nselect2 nselect2.n6 1.81877
R997 select0.n5 select0.t1 327.99
R998 select0.n9 select0.t5 293.969
R999 select0.n3 select0.t8 261.887
R1000 select0.n1 select0.t4 212.081
R1001 select0.n0 select0.t3 212.081
R1002 select0.n5 select0.t7 199.457
R1003 select0.n2 select0.n1 183.185
R1004 select0.n3 select0.t9 155.847
R1005 select0 select0.n9 154.065
R1006 select0.n6 select0.n5 152
R1007 select0.n4 select0.n3 152
R1008 select0.n1 select0.t2 139.78
R1009 select0.n0 select0.t0 139.78
R1010 select0.n9 select0.t6 138.338
R1011 select0.n1 select0.n0 61.346
R1012 select0.n10 select0 13.4199
R1013 select0.n8 select0.n4 11.9062
R1014 select0.n11 select0.n8 11.7395
R1015 select0.n12 select0.n11 11.5949
R1016 select0.n12 select0.n2 9.68118
R1017 select0.n7 select0 9.17383
R1018 select0.n2 select0 5.8885
R1019 select0.n10 select0 5.57469
R1020 select0.n8 select0.n7 4.6505
R1021 select0.n11 select0.n10 4.6505
R1022 select0.n7 select0.n6 2.98717
R1023 select0.n6 select0 2.34717
R1024 select0.n4 select0 2.07109
R1025 select0 select0.n12 0.559212
R1026 A2.n1 A2.t3 26.3998
R1027 A2.n1 A2.t2 23.5483
R1028 A2.n0 A2.t1 12.7127
R1029 A2.n0 A2.t0 10.8578
R1030 A2.n2 A2.n1 3.12177
R1031 A2.n2 A2.n0 1.81453
R1032 A2.n3 A2.n2 1.1255
R1033 A2.n3 A2 0.219402
R1034 A2 A2.n3 0.0655
R1035 A1.n1 A1.t0 26.3998
R1036 A1.n1 A1.t1 23.5483
R1037 A1.n0 A1.t3 12.7127
R1038 A1.n0 A1.t2 10.8578
R1039 A1.n2 A1.n1 3.12177
R1040 A1.n2 A1.n0 1.81453
R1041 A1.n3 A1.n2 1.1255
R1042 A1 A1.n3 0.21174
R1043 A1.n3 A1 0.0655
C0 m2_748_3404# mux4onehot_0.x2.GN1 0.06935f
C1 mux4onehot_0.x1.nSEL0 m2_748_3404# 3.43e-19
C2 A2 A1 1.81909f
C3 mux4onehot_0.select2 mux4onehot_0.x2.GN1 0.009187f
C4 select1 mux4onehot_0.x2.GN3 0.272312f
C5 mux4onehot_0.select2 mux4onehot_0.x1.nSEL0 0.131218f
C6 VDD nselect2 1.06761f
C7 a_617_4371# mux4onehot_0.x2.GN4 6.84e-19
C8 VDD mux4onehot_0.x1.nSEL1 0.481997f
C9 mux4onehot_0.x1.nSEL1 a_671_3541# 0.00175f
C10 select1 a_617_3819# 0.03417f
C11 A2 mux4onehot_0.x2.GN1 1.78e-19
C12 VDD Z 12.1648f
C13 mux4onehot_0.x2.GN4 m3_3538_4828# 7.17e-19
C14 VDD mux4onehot_0.x2.GP3 1.78265f
C15 a_617_4371# a_617_3995# 3.02e-19
C16 nselect2 a_617_4547# 6.01e-20
C17 A3 mux4onehot_0.x2.GN2 0.004147f
C18 mux4onehot_0.x2.GN2 a_617_5059# 7.58e-21
C19 mux4onehot_0.x1.nSEL1 a_617_4547# 1.59e-19
C20 a_643_4499# mux4onehot_0.x2.GN2 3.11e-20
C21 mux4onehot_0.x2.GN4 A4 3.83756f
C22 mux4onehot_0.x2.GN3 mux4onehot_0.x2.GN2 0.067582f
C23 select1 VDD 2.64545f
C24 mux4onehot_0.x2.GP3 a_617_4547# 5.21e-19
C25 a_617_3819# a_617_3403# 0.002207f
C26 mux4onehot_0.x2.GN2 a_617_3819# 0.106186f
C27 mux4onehot_0.x2.GN3 a_643_3947# 5.17e-20
C28 A2 mux4onehot_0.x2.GN4 3.42e-19
C29 mux4onehot_0.x2.GN4 m3_4582_4824# 7.07e-19
C30 mux4onehot_0.select2 a_617_3995# 1.67e-19
C31 mux4onehot_0.x2.GN3 A1 0.002069f
C32 m3_5612_4838# mux4onehot_0.x2.GP3 0.006132f
C33 a_617_3819# a_643_3947# 0.004764f
C34 select1 a_617_4547# 0.127717f
C35 mux4onehot_0.x2.GN3 mux4onehot_0.x2.GN1 0.002861f
C36 select0 nselect2 1.88e-19
C37 VDD a_617_3403# 0.210313f
C38 VDD mux4onehot_0.x2.GN2 0.60109f
C39 mux4onehot_0.x2.GN3 mux4onehot_0.x1.nSEL0 4.01e-20
C40 select0 mux4onehot_0.x1.nSEL1 0.168464f
C41 a_617_4371# mux4onehot_0.select2 0.009143f
C42 a_671_5197# a_617_5059# 0.006584f
C43 a_671_3541# a_617_3403# 0.006584f
C44 a_671_3541# mux4onehot_0.x2.GN2 8.86e-19
C45 a_617_3819# mux4onehot_0.x2.GN1 0.012466f
C46 select0 Z 4.1e-22
C47 mux4onehot_0.x1.nSEL0 a_617_3819# 0.03096f
C48 VDD a_643_3947# 4.32e-19
C49 mux4onehot_0.x2.GN3 a_671_5197# 1.07e-20
C50 select0 mux4onehot_0.x2.GP3 2.82e-19
C51 A3 mux4onehot_0.x2.GN4 0.187073f
C52 VDD A1 1.98654f
C53 mux4onehot_0.x2.GN2 a_617_4547# 5.62e-20
C54 mux4onehot_0.x2.GN4 a_617_5059# 0.134079f
C55 a_643_4499# mux4onehot_0.x2.GN4 3.22e-19
C56 mux4onehot_0.select2 m2_748_3404# 4.4e-19
C57 A2 m3_3538_4828# 0.1002f
C58 m3_4582_4824# m3_3538_4828# 0.003764f
C59 mux4onehot_0.x2.GN3 mux4onehot_0.x2.GN4 0.071502f
C60 VDD mux4onehot_0.x2.GN1 1.36577f
C61 select1 select0 1.66811f
C62 VDD mux4onehot_0.x1.nSEL0 0.391764f
C63 a_671_3541# mux4onehot_0.x2.GN1 0.001144f
C64 A1 a_617_4547# 5.02e-20
C65 A2 A4 2.39e-19
C66 m3_4582_4824# A4 6.07e-21
C67 mux4onehot_0.x2.GN3 a_617_3995# 0.048646f
C68 mux4onehot_0.x1.nSEL1 nselect2 0.047548f
C69 VDD a_671_5197# 8.97e-19
C70 a_617_4547# mux4onehot_0.x2.GN1 3.78e-20
C71 mux4onehot_0.x1.nSEL0 a_617_4547# 1.21e-20
C72 a_617_3819# a_617_3995# 0.185422f
C73 a_643_4499# a_617_4371# 0.004764f
C74 select0 a_617_3403# 0.048888f
C75 select0 mux4onehot_0.x2.GN2 0.114345f
C76 VDD mux4onehot_0.x2.GN4 1.23504f
C77 a_617_4371# mux4onehot_0.x2.GN3 0.104343f
C78 Z mux4onehot_0.x2.GP3 0.359536f
C79 select1 nselect2 0.001177f
C80 mux4onehot_0.x2.GN3 m3_3538_4828# 0.001446f
C81 VDD a_617_3995# 0.19314f
C82 select1 mux4onehot_0.x1.nSEL1 0.272823f
C83 select0 A1 3.49e-20
C84 A3 A4 2.08862f
C85 mux4onehot_0.x2.GN4 a_617_4547# 0.003699f
C86 select1 mux4onehot_0.x2.GP3 0.003386f
C87 mux4onehot_0.x2.GN3 A4 0.004656f
C88 select0 mux4onehot_0.x2.GN1 0.020307f
C89 mux4onehot_0.x2.GN3 mux4onehot_0.select2 0.001055f
C90 A3 A2 1.81997f
C91 select0 mux4onehot_0.x1.nSEL0 0.324538f
C92 m3_5612_4838# mux4onehot_0.x2.GN4 0.084813f
C93 A3 m3_4582_4824# 0.097296f
C94 a_617_4371# VDD 0.171441f
C95 mux4onehot_0.select2 a_617_3819# 8.66e-20
C96 mux4onehot_0.x2.GN3 A2 0.164396f
C97 select0 a_671_5197# 1.4e-19
C98 mux4onehot_0.x2.GN3 m3_4582_4824# 0.087318f
C99 mux4onehot_0.x1.nSEL1 a_617_3403# 0.193944f
C100 mux4onehot_0.x1.nSEL1 mux4onehot_0.x2.GN2 0.209956f
C101 Z mux4onehot_0.x2.GN2 0.429803f
C102 a_617_4371# a_617_4547# 0.185422f
C103 mux4onehot_0.x1.nSEL1 a_643_3947# 9.57e-19
C104 mux4onehot_0.x2.GN2 mux4onehot_0.x2.GP3 0.004319f
C105 VDD m2_748_3404# 0.139545f
C106 select0 mux4onehot_0.x2.GN4 0.218396f
C107 VDD A4 1.54289f
C108 VDD mux4onehot_0.select2 0.231538f
C109 Z A1 4.52f
C110 select1 a_617_3403# 0.02803f
C111 A1 mux4onehot_0.x2.GP3 0.001277f
C112 select0 a_617_3995# 0.143958f
C113 select1 mux4onehot_0.x2.GN2 0.108649f
C114 mux4onehot_0.x1.nSEL1 mux4onehot_0.x2.GN1 0.034891f
C115 VDD A2 1.61513f
C116 mux4onehot_0.x1.nSEL1 mux4onehot_0.x1.nSEL0 0.352716f
C117 Z mux4onehot_0.x2.GN1 0.428922f
C118 mux4onehot_0.x2.GN3 A3 3.80503f
C119 mux4onehot_0.x2.GN3 a_617_5059# 1.07e-20
C120 mux4onehot_0.x2.GP3 mux4onehot_0.x2.GN1 0.002439f
C121 a_643_4499# mux4onehot_0.x2.GN3 0.001073f
C122 select1 A1 1.45e-21
C123 m3_5612_4838# A4 0.091998f
C124 a_617_4371# select0 0.086353f
C125 mux4onehot_0.x2.GN3 a_617_3819# 6.68e-19
C126 select1 mux4onehot_0.x2.GN1 0.312198f
C127 mux4onehot_0.x2.GN4 nselect2 1.53e-20
C128 mux4onehot_0.x2.GN2 a_617_3403# 0.039612f
C129 select1 mux4onehot_0.x1.nSEL0 0.137403f
C130 m3_5612_4838# m3_4582_4824# 0.003741f
C131 Z mux4onehot_0.x2.GN4 0.44705f
C132 VDD A3 1.61205f
C133 mux4onehot_0.x2.GN2 a_643_3947# 0.002418f
C134 VDD a_617_5059# 0.217381f
C135 select0 m2_748_3404# 0.130999f
C136 mux4onehot_0.x2.GP3 mux4onehot_0.x2.GN4 3.44338f
C137 select1 a_671_5197# 8.84e-19
C138 a_643_4499# VDD 0.001496f
C139 mux4onehot_0.x1.nSEL1 a_617_3995# 0.041068f
C140 mux4onehot_0.x2.GN2 A1 0.157008f
C141 select0 mux4onehot_0.select2 0.368835f
C142 VDD mux4onehot_0.x2.GN3 0.650424f
C143 a_617_3403# mux4onehot_0.x2.GN1 0.12869f
C144 mux4onehot_0.x2.GN2 mux4onehot_0.x2.GN1 0.065209f
C145 VDD a_617_3819# 0.161854f
C146 select1 mux4onehot_0.x2.GN4 0.059813f
C147 mux4onehot_0.x1.nSEL0 a_617_3403# 0.081627f
C148 mux4onehot_0.x1.nSEL0 mux4onehot_0.x2.GN2 0.154394f
C149 a_617_4371# nselect2 1.29e-19
C150 a_617_4371# mux4onehot_0.x1.nSEL1 7.84e-19
C151 mux4onehot_0.x2.GN3 a_617_4547# 0.004288f
C152 a_643_3947# mux4onehot_0.x2.GN1 1.22e-20
C153 mux4onehot_0.x1.nSEL0 a_643_3947# 2.51e-19
C154 a_671_5197# mux4onehot_0.x2.GN2 8.14e-21
C155 select1 a_617_3995# 0.254026f
C156 A1 mux4onehot_0.x2.GN1 4.61829f
C157 a_617_4371# mux4onehot_0.x2.GP3 0.00144f
C158 mux4onehot_0.x1.nSEL0 A1 1.93e-21
C159 m3_5612_4838# mux4onehot_0.x2.GN3 0.016026f
C160 VDD a_671_3541# 9.09e-19
C161 mux4onehot_0.x1.nSEL1 m2_748_3404# 0.00815f
C162 mux4onehot_0.x2.GP3 m3_3538_4828# 9.67e-19
C163 mux4onehot_0.x2.GN2 mux4onehot_0.x2.GN4 8.84e-19
C164 mux4onehot_0.select2 nselect2 0.150826f
C165 mux4onehot_0.x1.nSEL0 mux4onehot_0.x2.GN1 0.004383f
C166 mux4onehot_0.select2 mux4onehot_0.x1.nSEL1 0.164723f
C167 select1 a_617_4371# 0.261734f
C168 Z A4 4.51511f
C169 VDD a_617_4547# 0.262185f
C170 select0 a_617_5059# 0.220366f
C171 mux4onehot_0.x2.GP3 A4 0.161499f
C172 a_643_4499# select0 0.001558f
C173 mux4onehot_0.x2.GN2 a_617_3995# 0.017018f
C174 A1 mux4onehot_0.x2.GN4 0.001437f
C175 select0 mux4onehot_0.x2.GN3 0.254198f
C176 Z A2 4.52054f
C177 select1 m2_748_3404# 0.183786f
C178 A2 mux4onehot_0.x2.GP3 0.001826f
C179 select0 a_617_3819# 0.246189f
C180 mux4onehot_0.x2.GN4 mux4onehot_0.x2.GN1 0.001075f
C181 mux4onehot_0.x2.GP3 m3_4582_4824# 0.002824f
C182 select1 mux4onehot_0.select2 0.139336f
C183 mux4onehot_0.x1.nSEL0 mux4onehot_0.x2.GN4 2.26e-20
C184 a_617_4371# mux4onehot_0.x2.GN2 1.63e-19
C185 a_617_3995# mux4onehot_0.x2.GN1 1.46e-19
C186 a_671_5197# mux4onehot_0.x2.GN4 0.001562f
C187 mux4onehot_0.x2.GN2 m3_3538_4828# 0.099332f
C188 mux4onehot_0.x1.nSEL0 a_617_3995# 0.001174f
C189 select0 VDD 1.09594f
C190 a_617_4371# A1 1.55e-21
C191 nselect2 a_617_5059# 9.77e-20
C192 select0 a_671_3541# 9.55e-19
C193 a_617_3403# m2_748_3404# 0.01297f
C194 a_643_4499# mux4onehot_0.x1.nSEL1 4.08e-19
C195 Z A3 4.52142f
C196 mux4onehot_0.select2 mux4onehot_0.x2.GN2 0.001308f
C197 mux4onehot_0.x2.GN3 nselect2 7.39e-21
C198 a_617_4371# mux4onehot_0.x2.GN1 6.43e-20
C199 mux4onehot_0.x2.GN3 mux4onehot_0.x1.nSEL1 0.012418f
C200 A3 mux4onehot_0.x2.GP3 4.01143f
C201 a_617_4371# mux4onehot_0.x1.nSEL0 1.91e-20
C202 select0 a_617_4547# 0.279858f
C203 a_643_4499# mux4onehot_0.x2.GP3 4.39e-19
C204 mux4onehot_0.x2.GN3 Z 0.4304f
C205 mux4onehot_0.x1.nSEL1 a_617_3819# 0.073392f
C206 mux4onehot_0.x2.GN2 A2 3.81462f
C207 m3_3538_4828# mux4onehot_0.x2.GN1 6.03e-20
C208 mux4onehot_0.x2.GN2 m3_4582_4824# 0.016745f
C209 mux4onehot_0.x2.GN3 mux4onehot_0.x2.GP3 2.87029f
C210 select1 a_617_5059# 0.125445f
C211 A4 VSS 3.673693f
C212 A3 VSS 3.139098f
C213 A2 VSS 3.238408f
C214 Z VSS 13.09264f
C215 A1 VSS 3.972022f
C216 nselect2 VSS 0.47102f
C217 select0 VSS 1.41757f
C218 select1 VSS 1.610707f
C219 VDD VSS 55.994358f
C220 m3_5612_4838# VSS 0.090191f $ **FLOATING
C221 m3_4582_4824# VSS 0.086003f $ **FLOATING
C222 m3_3538_4828# VSS 0.168273f $ **FLOATING
C223 m2_748_3404# VSS 0.065655f $ **FLOATING
C224 a_671_3541# VSS 0.006505f
C225 a_617_3403# VSS 0.266782f
C226 mux4onehot_0.x1.nSEL0 VSS 0.649982f
C227 mux4onehot_0.x2.GN1 VSS 6.356356f
C228 a_643_3947# VSS 0.004461f
C229 a_617_3819# VSS 0.220868f
C230 mux4onehot_0.x1.nSEL1 VSS 0.69132f
C231 mux4onehot_0.x2.GN2 VSS 3.93113f
C232 a_617_3995# VSS 0.23458f
C233 mux4onehot_0.select2 VSS 1.16504f
C234 mux4onehot_0.x2.GP3 VSS 1.67016f
C235 a_643_4499# VSS 0.006801f
C236 mux4onehot_0.x2.GN3 VSS 3.6536f
C237 a_617_4371# VSS 0.232764f
C238 a_617_4547# VSS 0.249604f
C239 mux4onehot_0.x2.GN4 VSS 7.589221f
C240 a_671_5197# VSS 0.006439f
C241 a_617_5059# VSS 0.306675f
C242 A1.t3 VSS 0.813767f
C243 A1.t2 VSS 0.467169f
C244 A1.n0 VSS 4.5246f
C245 A1.t0 VSS 0.842259f
C246 A1.t1 VSS 0.59582f
C247 A1.n1 VSS 4.62603f
C248 A1.n2 VSS 0.731719f
C249 A1.n3 VSS 0.224671f
C250 A2.t1 VSS 0.763965f
C251 A2.t0 VSS 0.438578f
C252 A2.n0 VSS 4.2477f
C253 A2.t3 VSS 0.790712f
C254 A2.t2 VSS 0.559356f
C255 A2.n1 VSS 4.34292f
C256 A2.n2 VSS 0.686937f
C257 A2.n3 VSS 0.222065f
C258 mux4onehot_0.x2.GN4.t0 VSS 0.060733f
C259 mux4onehot_0.x2.GN4.n0 VSS 0.070011f
C260 mux4onehot_0.x2.GN4.t6 VSS 0.686349f
C261 mux4onehot_0.x2.GN4.t4 VSS 0.66979f
C262 mux4onehot_0.x2.GN4.n1 VSS 3.00509f
C263 mux4onehot_0.x2.GN4.n2 VSS 1.54925f
C264 mux4onehot_0.x2.GN4.t3 VSS 0.038126f
C265 mux4onehot_0.x2.GN4.t7 VSS 0.022467f
C266 mux4onehot_0.x2.GN4.t2 VSS 0.038126f
C267 mux4onehot_0.x2.GN4.t5 VSS 0.022467f
C268 mux4onehot_0.x2.GN4.n3 VSS 0.06397f
C269 mux4onehot_0.x2.GN4.n4 VSS 0.094764f
C270 mux4onehot_0.x2.GN4.n5 VSS 0.042424f
C271 mux4onehot_0.x2.GN4.n6 VSS 0.343642f
C272 mux4onehot_0.x2.GN4.t1 VSS 0.155108f
C273 mux4onehot_0.x2.GN4.n7 VSS 0.027899f
C274 mux4onehot_0.x2.GN4.n8 VSS 0.031254f
C275 A4.t3 VSS 0.893325f
C276 A4.t0 VSS 0.512841f
C277 A4.n0 VSS 4.96695f
C278 A4.t1 VSS 0.924602f
C279 A4.t2 VSS 0.65407f
C280 A4.n1 VSS 5.0783f
C281 A4.n2 VSS 0.803255f
C282 A4.n3 VSS 0.258761f
C283 mux4onehot_0.x2.GP4.n0 VSS 0.095571f
C284 mux4onehot_0.x2.x4.GP VSS 2.50543f
C285 mux4onehot_0.x1.gpo3 VSS 1.18077f
C286 mux4onehot_0.x2.GP4.t1 VSS 0.012052f
C287 mux4onehot_0.x2.GP4.t0 VSS 0.012052f
C288 mux4onehot_0.x2.GP4.n1 VSS 0.028739f
C289 mux4onehot_0.x1.x14.Y VSS 0.104168f
C290 mux4onehot_0.x2.GP4.t4 VSS 0.609957f
C291 mux4onehot_0.x2.GP4.t5 VSS 0.626965f
C292 mux4onehot_0.x2.GP4.n2 VSS 2.22891f
C293 mux4onehot_0.x2.GP4.n3 VSS 0.017567f
C294 mux4onehot_0.x2.GP4.t2 VSS 0.018542f
C295 mux4onehot_0.x2.GP4.t3 VSS 0.018542f
C296 mux4onehot_0.x2.GP4.n4 VSS 0.040723f
C297 select1.t6 VSS 0.032343f
C298 select1.t4 VSS 0.019059f
C299 select1.t3 VSS 0.032343f
C300 select1.t2 VSS 0.019059f
C301 select1.n0 VSS 0.054267f
C302 select1.n1 VSS 0.080179f
C303 select1.n2 VSS 0.048819f
C304 select1.t9 VSS 0.014966f
C305 select1.t0 VSS 0.031563f
C306 select1.n3 VSS 0.113336f
C307 select1.n4 VSS 0.021975f
C308 select1.n5 VSS 0.018928f
C309 select1.t5 VSS 0.022802f
C310 select1.t7 VSS 0.015669f
C311 select1.n6 VSS 0.06626f
C312 select1.n7 VSS 0.015263f
C313 select1.n8 VSS 0.109332f
C314 select1.n9 VSS 0.396f
C315 select1.t8 VSS 0.02778f
C316 select1.t1 VSS 0.018863f
C317 select1.n10 VSS 0.065634f
C318 select1.n11 VSS 0.01571f
C319 select1.n12 VSS 0.101902f
C320 select1.n13 VSS 0.457083f
C321 select1.n14 VSS 0.597136f
C322 mux4onehot_0.x2.x2.GP VSS 2.76866f
C323 mux4onehot_0.x1.gpo1 VSS 0.998586f
C324 mux4onehot_0.x2.GP2.t1 VSS 0.016016f
C325 mux4onehot_0.x2.GP2.t0 VSS 0.016016f
C326 mux4onehot_0.x2.GP2.n0 VSS 0.03819f
C327 mux4onehot_0.x1.x12.Y VSS 0.058128f
C328 mux4onehot_0.x2.GP2.n1 VSS 0.075027f
C329 mux4onehot_0.x2.GP2.n2 VSS 0.023344f
C330 mux4onehot_0.x2.GP2.t3 VSS 0.02464f
C331 mux4onehot_0.x2.GP2.t2 VSS 0.02464f
C332 mux4onehot_0.x2.GP2.n3 VSS 0.050813f
C333 mux4onehot_0.x2.GP2.t5 VSS 0.810542f
C334 mux4onehot_0.x2.GP2.t4 VSS 0.833144f
C335 mux4onehot_0.x2.GP2.n4 VSS 2.95587f
C336 mux4onehot_0.x2.GP2.n5 VSS 0.106388f
C337 Z.t6 VSS 0.331048f
C338 Z.n0 VSS 0.494313f
C339 Z.t5 VSS 0.337693f
C340 Z.t4 VSS 0.448126f
C341 Z.n1 VSS 2.26138f
C342 Z.n2 VSS 0.765155f
C343 Z.t3 VSS 0.436117f
C344 Z.n3 VSS 0.542399f
C345 Z.n4 VSS 0.689241f
C346 Z.t8 VSS 0.331048f
C347 Z.n5 VSS 0.494313f
C348 Z.t7 VSS 0.337693f
C349 Z.t0 VSS 0.448126f
C350 Z.n6 VSS 2.26138f
C351 Z.n7 VSS 0.765155f
C352 Z.t14 VSS 0.436117f
C353 Z.n8 VSS 0.542399f
C354 Z.n9 VSS 0.668421f
C355 Z.n10 VSS 0.295408f
C356 Z.t13 VSS 0.331048f
C357 Z.n11 VSS 0.494313f
C358 Z.t12 VSS 0.337693f
C359 Z.t11 VSS 0.448126f
C360 Z.n12 VSS 2.26138f
C361 Z.n13 VSS 0.765155f
C362 Z.t10 VSS 0.436117f
C363 Z.n14 VSS 0.542399f
C364 Z.n15 VSS 0.666353f
C365 Z.n16 VSS 0.303503f
C366 Z.t15 VSS 0.331048f
C367 Z.n17 VSS 0.494313f
C368 Z.t9 VSS 0.337693f
C369 Z.t1 VSS 0.448126f
C370 Z.n18 VSS 2.26138f
C371 Z.n19 VSS 0.765155f
C372 Z.t2 VSS 0.436117f
C373 Z.n20 VSS 0.542399f
C374 Z.n21 VSS 0.679854f
C375 Z.n22 VSS 0.354074f
C376 Z.n23 VSS 0.796049f
C377 Z.n24 VSS 0.726738f
C378 A3.t2 VSS 0.893857f
C379 A3.t3 VSS 0.513146f
C380 A3.n0 VSS 4.9699f
C381 A3.t1 VSS 0.925152f
C382 A3.t0 VSS 0.654459f
C383 A3.n1 VSS 5.08132f
C384 A3.n2 VSS 0.803733f
C385 A3.n3 VSS 0.264783f
C386 VDD.n0 VSS 0.004385f
C387 VDD.t36 VSS 0.008849f
C388 VDD.n1 VSS 0.008705f
C389 VDD.t58 VSS 9.5e-19
C390 VDD.t40 VSS 0.001443f
C391 VDD.n2 VSS 0.002493f
C392 VDD.t34 VSS 0.00902f
C393 VDD.t32 VSS 0.008849f
C394 VDD.n3 VSS 0.008429f
C395 VDD.n4 VSS 0.004385f
C396 VDD.n5 VSS 0.003969f
C397 VDD.t20 VSS 0.001302f
C398 VDD.n6 VSS 0.003696f
C399 VDD.t38 VSS 0.005354f
C400 VDD.n7 VSS 0.004928f
C401 VDD.n8 VSS 0.004398f
C402 VDD.t30 VSS 0.008852f
C403 VDD.n9 VSS 7.24e-19
C404 VDD.t27 VSS 0.003795f
C405 VDD.t13 VSS 0.006265f
C406 VDD.n10 VSS 0.006176f
C407 VDD.n11 VSS 0.007402f
C408 VDD.t71 VSS 0.026146f
C409 VDD.n12 VSS 0.023649f
C410 VDD.t56 VSS 7.09e-19
C411 VDD.t50 VSS 0.001902f
C412 VDD.n13 VSS 0.00868f
C413 VDD.t14 VSS 0.006265f
C414 VDD.n14 VSS 0.004584f
C415 VDD.n15 VSS 0.017109f
C416 VDD.n16 VSS 0.013517f
C417 VDD.n17 VSS 0.017558f
C418 VDD.n18 VSS 0.010138f
C419 VDD.n19 VSS 0.007402f
C420 VDD.n20 VSS 0.005552f
C421 VDD.n21 VSS 0.003485f
C422 VDD.n22 VSS 0.010979f
C423 VDD.n23 VSS 0.017211f
C424 VDD.t45 VSS 0.017789f
C425 VDD.n24 VSS 0.001339f
C426 VDD.n25 VSS 0.001368f
C427 VDD.n26 VSS 0.005552f
C428 VDD.n27 VSS 0.00171f
C429 VDD.t60 VSS 0.008971f
C430 VDD.n28 VSS 0.007362f
C431 VDD.n29 VSS 0.004385f
C432 VDD.t72 VSS 0.026146f
C433 VDD.n30 VSS 0.006517f
C434 VDD.n31 VSS 0.004385f
C435 VDD.t62 VSS 7.09e-19
C436 VDD.t66 VSS 0.001902f
C437 VDD.n32 VSS 0.00868f
C438 VDD.t73 VSS 0.026146f
C439 VDD.t64 VSS 0.003795f
C440 VDD.n33 VSS 0.01172f
C441 VDD.n34 VSS 0.006718f
C442 VDD.n35 VSS 0.003485f
C443 VDD.t4 VSS 0.006265f
C444 VDD.n36 VSS 0.006176f
C445 VDD.n37 VSS 0.023649f
C446 VDD.n38 VSS 0.010138f
C447 VDD.n39 VSS 0.017558f
C448 VDD.t5 VSS 0.006265f
C449 VDD.t23 VSS 0.008972f
C450 VDD.n40 VSS 0.002534f
C451 VDD.n41 VSS 0.003017f
C452 VDD.t63 VSS 0.035816f
C453 VDD.t65 VSS 0.03463f
C454 VDD.t3 VSS 0.025617f
C455 VDD.t61 VSS 0.036764f
C456 VDD.t53 VSS 0.035816f
C457 VDD.t1 VSS 0.040797f
C458 VDD.t47 VSS 0.029649f
C459 VDD.t24 VSS 0.015892f
C460 VDD.t59 VSS 0.007353f
C461 VDD.t22 VSS 0.025854f
C462 VDD.n42 VSS 0.033737f
C463 VDD.n43 VSS 0.023396f
C464 VDD.n44 VSS 0.006877f
C465 VDD.n45 VSS 0.011034f
C466 VDD.n46 VSS 0.013517f
C467 VDD.n47 VSS 0.004586f
C468 VDD.n48 VSS 0.036532f
C469 VDD.n49 VSS 0.049693f
C470 VDD.t10 VSS 0.006265f
C471 VDD.n50 VSS 0.012251f
C472 VDD.n51 VSS 0.023649f
C473 VDD.n52 VSS 0.014573f
C474 VDD.t11 VSS 0.006265f
C475 VDD.t42 VSS 0.009015f
C476 VDD.n53 VSS 0.010534f
C477 VDD.t9 VSS 0.080577f
C478 VDD.t6 VSS 0.049502f
C479 VDD.t17 VSS 0.020312f
C480 VDD.t67 VSS 0.028114f
C481 VDD.t69 VSS 0.020312f
C482 VDD.t15 VSS 0.028114f
C483 VDD.t43 VSS 0.020312f
C484 VDD.t41 VSS 0.030401f
C485 VDD.n54 VSS 0.033279f
C486 VDD.n55 VSS 0.004385f
C487 VDD.n56 VSS 0.001909f
C488 VDD.t16 VSS 0.009015f
C489 VDD.n57 VSS 0.001909f
C490 VDD.t68 VSS 0.009015f
C491 VDD.n58 VSS 0.128854f
C492 VDD.n59 VSS 0.007542f
C493 VDD.n60 VSS 0.004584f
C494 VDD.t74 VSS 0.026555f
C495 VDD.t7 VSS 0.006265f
C496 VDD.n61 VSS 0.026289f
C497 VDD.n62 VSS 0.013065f
C498 VDD.t8 VSS 0.006265f
C499 VDD.n63 VSS 0.017109f
C500 VDD.n64 VSS 0.015735f
C501 VDD.n65 VSS 0.009873f
C502 VDD.n66 VSS 0.007705f
C503 VDD.n67 VSS 0.007513f
C504 VDD.t18 VSS 0.00902f
C505 VDD.n68 VSS 0.011351f
C506 VDD.n69 VSS 0.004385f
C507 VDD.n70 VSS 0.007402f
C508 VDD.n71 VSS 0.005552f
C509 VDD.n72 VSS 0.010648f
C510 VDD.t70 VSS 0.00902f
C511 VDD.n73 VSS 0.011522f
C512 VDD.n74 VSS 0.004385f
C513 VDD.n75 VSS 0.007402f
C514 VDD.n76 VSS 0.005552f
C515 VDD.n77 VSS 0.010648f
C516 VDD.t44 VSS 0.00902f
C517 VDD.n78 VSS 0.011522f
C518 VDD.n79 VSS 0.001909f
C519 VDD.n80 VSS 0.007402f
C520 VDD.n81 VSS 0.005552f
C521 VDD.n82 VSS 0.002816f
C522 VDD.n83 VSS 0.015383f
C523 VDD.n84 VSS 0.006877f
C524 VDD.n85 VSS 0.011034f
C525 VDD.n86 VSS 0.018798f
C526 VDD.n87 VSS 0.003741f
C527 VDD.n88 VSS 0.033997f
C528 VDD.n89 VSS 0.032966f
C529 VDD.n90 VSS 7.64e-19
C530 VDD.t25 VSS 9.5e-19
C531 VDD.t48 VSS 0.001443f
C532 VDD.n91 VSS 0.002493f
C533 VDD.n92 VSS 0.016734f
C534 VDD.t52 VSS 0.009015f
C535 VDD.n93 VSS 0.010506f
C536 VDD.t2 VSS 0.00297f
C537 VDD.t46 VSS 0.007895f
C538 VDD.n94 VSS 0.004479f
C539 VDD.t54 VSS 0.008852f
C540 VDD.n95 VSS 0.009339f
C541 VDD.n96 VSS 0.012012f
C542 VDD.n97 VSS 0.001582f
C543 VDD.n98 VSS 0.007402f
C544 VDD.n99 VSS 0.004385f
C545 VDD.n100 VSS 0.002534f
C546 VDD.n101 VSS 0.002816f
C547 VDD.n102 VSS 0.015073f
C548 VDD.n103 VSS 0.041101f
C549 VDD.t57 VSS 0.007827f
C550 VDD.t35 VSS 0.020398f
C551 VDD.t33 VSS 0.02277f
C552 VDD.t39 VSS 0.015892f
C553 VDD.t19 VSS 0.029649f
C554 VDD.t31 VSS 0.041745f
C555 VDD.t29 VSS 0.020398f
C556 VDD.t37 VSS 0.015892f
C557 VDD.t55 VSS 0.036764f
C558 VDD.t12 VSS 0.025617f
C559 VDD.t49 VSS 0.03463f
C560 VDD.t26 VSS 0.035816f
C561 VDD.n104 VSS 0.02439f
C562 VDD.n105 VSS 0.007086f
C563 VDD.n106 VSS 0.005044f
C564 VDD.n107 VSS 0.001339f
C565 VDD.n108 VSS 0.009827f
C566 VDD.n109 VSS 0.003748f
C567 VDD.n110 VSS 0.007402f
C568 VDD.n111 VSS 0.005552f
C569 VDD.n112 VSS 0.0033f
C570 VDD.n113 VSS 0.011218f
C571 VDD.n114 VSS 0.008028f
C572 VDD.n115 VSS 0.005109f
C573 VDD.n116 VSS 0.014448f
C574 VDD.n117 VSS 0.091894f
C575 VDD.n118 VSS 0.196687f
C576 VDD.n119 VSS 0.258918f
C577 VDD.n120 VSS 0.143929f
C578 VDD.n121 VSS 0.032339f
C579 VDD.n122 VSS 0.143929f
C580 VDD.n123 VSS 0.069513f
C581 VDD.n124 VSS 0.585446f
C582 VDD.n125 VSS 0.585446f
C583 VDD.n126 VSS 0.096355f
C584 VDD.n127 VSS 0.070572f
C585 VDD.t21 VSS 0.778437f
C586 VDD.n130 VSS 0.070572f
C587 VDD.n131 VSS 2.99e-19
C588 VDD.n132 VSS 0.042855f
C589 VDD.n133 VSS 0.007792f
C590 VDD.n134 VSS 0.084714f
C591 VDD.n135 VSS 0.045296f
C592 VDD.n136 VSS 0.09198f
C593 VDD.n137 VSS 0.106709f
C594 VDD.n138 VSS 0.143929f
C595 VDD.n139 VSS 0.002337f
C596 VDD.n140 VSS 0.096355f
C597 VDD.n141 VSS 0.070572f
C598 VDD.t51 VSS 0.778437f
C599 VDD.n143 VSS 0.585446f
C600 VDD.n144 VSS 0.070572f
C601 VDD.n146 VSS 0.585446f
C602 VDD.n147 VSS 0.069513f
C603 VDD.n148 VSS 0.005595f
C604 VDD.n149 VSS 0.042812f
C605 VDD.n150 VSS 0.007863f
C606 VDD.n151 VSS 0.084714f
C607 VDD.n152 VSS 0.044937f
C608 VDD.n153 VSS 0.072829f
C609 VDD.n154 VSS 0.104614f
C610 VDD.n155 VSS 0.143929f
C611 VDD.n156 VSS 0.002479f
C612 VDD.n157 VSS 0.096355f
C613 VDD.n158 VSS 0.070572f
C614 VDD.t0 VSS 0.778437f
C615 VDD.n160 VSS 0.585446f
C616 VDD.n161 VSS 0.070572f
C617 VDD.n163 VSS 0.585446f
C618 VDD.n164 VSS 0.069513f
C619 VDD.n165 VSS 0.005604f
C620 VDD.n166 VSS 0.042669f
C621 VDD.n167 VSS 0.007863f
C622 VDD.n168 VSS 0.084714f
C623 VDD.n169 VSS 0.044937f
C624 VDD.n170 VSS 0.070999f
C625 VDD.n171 VSS 0.108876f
C626 VDD.n172 VSS 0.007654f
C627 VDD.n173 VSS 0.069513f
C628 VDD.n174 VSS 0.585446f
C629 VDD.n175 VSS 0.585446f
C630 VDD.n176 VSS 0.096355f
C631 VDD.n177 VSS 0.070572f
C632 VDD.t28 VSS 0.778437f
C633 VDD.n180 VSS 0.070572f
C634 VDD.n181 VSS 2.71e-19
C635 VDD.n182 VSS 0.042855f
C636 VDD.n183 VSS 0.007821f
C637 VDD.n184 VSS 0.084714f
C638 VDD.n185 VSS 0.045267f
C639 mux4onehot_0.x2.x1.GP VSS 1.98566f
C640 mux4onehot_0.x2.GP1.t2 VSS 0.012716f
C641 mux4onehot_0.x2.GP1.t3 VSS 0.012716f
C642 mux4onehot_0.x2.GP1.n0 VSS 0.03032f
C643 mux4onehot_0.x1.x11.Y VSS 0.046385f
C644 mux4onehot_0.x2.GP1.n1 VSS 0.059566f
C645 mux4onehot_0.x2.GP1.n2 VSS 0.018534f
C646 mux4onehot_0.x2.GP1.t0 VSS 0.019563f
C647 mux4onehot_0.x2.GP1.t1 VSS 0.019563f
C648 mux4onehot_0.x2.GP1.n3 VSS 0.040309f
C649 mux4onehot_0.x2.GP1.t4 VSS 0.643518f
C650 mux4onehot_0.x2.GP1.t5 VSS 0.661463f
C651 mux4onehot_0.x2.GP1.n4 VSS 2.33672f
C652 mux4onehot_0.x1.gpo0 VSS 0.626909f
C653 mux4onehot_0.x2.GP1.n5 VSS 0.086057f
C654 mux4onehot_0.x2.GN1.t0 VSS 0.029982f
C655 mux4onehot_0.x2.GN1.n0 VSS 0.034597f
C656 mux4onehot_0.x2.GN1.t5 VSS 0.338823f
C657 mux4onehot_0.x2.GN1.t7 VSS 0.330648f
C658 mux4onehot_0.x2.GN1.n1 VSS 1.48349f
C659 mux4onehot_0.x2.GN1.n2 VSS 0.518161f
C660 mux4onehot_0.x2.GN1.t6 VSS 0.018821f
C661 mux4onehot_0.x2.GN1.t3 VSS 0.011091f
C662 mux4onehot_0.x2.GN1.t4 VSS 0.018821f
C663 mux4onehot_0.x2.GN1.t2 VSS 0.011091f
C664 mux4onehot_0.x2.GN1.n3 VSS 0.031579f
C665 mux4onehot_0.x2.GN1.n4 VSS 0.046643f
C666 mux4onehot_0.x2.GN1.n5 VSS 0.045366f
C667 mux4onehot_0.x2.GN1.n6 VSS 0.098537f
C668 mux4onehot_0.x2.GN1.t1 VSS 0.076571f
C669 mux4onehot_0.x2.GN1.n7 VSS 0.013773f
C670 mux4onehot_0.x2.GN1.n8 VSS 0.015429f
.ends

