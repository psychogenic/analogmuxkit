** sch_path: /home/ttuser/vmswap/analogmuxkit/xschem/tb_mux8to1.sch
**.subckt tb_mux8to1
V2 net1 VSS sin(0.9 0.9 250k)
V3 net2 VSS sin(0.9 0.9 5Meg)
V5 net3 VSS sin(0.9 0.9 500k)
V6 net4 VSS sin(0.9 0.9 1Meg)
R2 IN1 net1 1 m=1
R3 IN2 net3 1 m=1
R4 IN3 net4 1 m=1
R5 IN4 net2 1 m=1
x1 SEL1 SEL2 IN1 IN3 IN2 IN4 OUT IN8 SEL0 IN7 IN6 VCC IN5 VSS mux8to1_parax
V1 net5 VSS dc 0.25 sin(0.3 0.1 1Meg)
R1 IN5 net5 1 m=1
V4 net6 VSS dc 0.88 sin(0.6 0.3 500k)
R6 IN6 net6 1 m=1
V7 net7 VSS dc 1.25
R7 IN7 net7 1 m=1
V8 net8 VSS dc 1.2 sin(1.2 0.4 200k)
R8 IN8 net8 1 m=1
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ttuser/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  mux8to1.sym # of pins=14
** sym_path: /home/ttuser/vmswap/analogmuxkit/xschem/mux8to1.sym
** sch_path: /home/ttuser/vmswap/analogmuxkit/xschem/mux8to1.sch
.subckt mux8to1 select0 select1 select2 A1 A2 A3 A4 A5 A6 A7 A8 Z VDD VSS
*.ipin select0
*.ipin select1
*.ipin select2
*.ipin VDD
*.ipin VSS
*.iopin Z
*.iopin A1
*.iopin A2
*.iopin A3
*.iopin A4
*.iopin A5
*.iopin A6
*.iopin A7
*.iopin A8
x4 OUT_HIGH select2 nSEL2 Z VDD VSS passgate
x5 OUT_LOW nSEL2 select2 Z VDD VSS passgate
x2 A1 gno0 gpo0 OUT_LOW A2 gno1 gpo1 OUT_LOW A3 gno2 gpo2 OUT_LOW A4 gno3 gpo3 OUT_LOW VDD VSS passgatex4
x1 select0 select1 select2 gno0 gpo0 gno1 gpo1 gno2 gpo2 gno3 gpo3 nSEL2 VDD VSS passgatesCtrlManual
x3 A5 gno0 gpo0 OUT_HIGH A6 gno1 gpo1 OUT_HIGH A7 gno2 gpo2 OUT_HIGH A8 gno3 gpo3 OUT_HIGH VDD VSS passgatex4
.ends


* expanding   symbol:  mux8to1_parax.sym # of pins=14
** sym_path: /home/ttuser/vmswap/analogmuxkit/xschem/mux8to1.sym
.include /home/ttuser/vmswap/analogmuxkit/xschem/extracted/mux8to1_parax.spice

* expanding   symbol:  passgate.sym # of pins=6
** sym_path: /home/ttuser/vmswap/analogmuxkit/xschem/passgate.sym
** sch_path: /home/ttuser/vmswap/analogmuxkit/xschem/passgate.sch
.subckt passgate A GN GP Z VDD VSS
*.ipin GN
*.ipin VDD
*.ipin VSS
*.ipin GP
*.iopin A
*.iopin Z
XM1 Z GN A VSS sky130_fd_pr__nfet_01v8_lvt L=0.35 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
XM3 Z GP A VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=2 m=2
.ends


* expanding   symbol:  passgatex4.sym # of pins=18
** sym_path: /home/ttuser/vmswap/analogmuxkit/xschem/passgatex4.sym
** sch_path: /home/ttuser/vmswap/analogmuxkit/xschem/passgatex4.sch
.subckt passgatex4 A1 GN1 GP1 Z1 A2 GN2 GP2 Z2 A3 GN3 GP3 Z3 A4 GN4 GP4 Z4 VDD VSS
*.ipin VDD
*.ipin VSS
*.ipin GP1
*.ipin GN1
*.iopin A1
*.iopin Z1
*.ipin GP2
*.ipin GN2
*.iopin A2
*.iopin Z2
*.ipin GP3
*.ipin GN3
*.iopin A3
*.iopin Z3
*.ipin GP4
*.ipin GN4
*.iopin A4
*.iopin Z4
x1 A1 GN1 GP1 Z1 VDD VSS passgate
x2 A2 GN2 GP2 Z2 VDD VSS passgate
x3 A3 GN3 GP3 Z3 VDD VSS passgate
x4 A4 GN4 GP4 Z4 VDD VSS passgate
.ends


* expanding   symbol:  passgatesCtrlManual.sym # of pins=14
** sym_path: /home/ttuser/vmswap/analogmuxkit/xschem/passgatesCtrlManual.sym
** sch_path: /home/ttuser/vmswap/analogmuxkit/xschem/passgatesCtrlManual.sch
.subckt passgatesCtrlManual SEL0 SEL1 SEL2 gno0 gpo0 gno1 gpo1 gno2 gpo2 gno3 gpo3 nSEL2 VPWR VGND
*.ipin SEL0
*.ipin SEL1
*.ipin SEL2
*.opin gno0
*.opin gpo0
*.opin gno1
*.opin gpo1
*.opin gno2
*.opin gpo2
*.opin gno3
*.opin gpo3
*.opin nSEL2
*.ipin VPWR
*.ipin VGND
x1 SEL0 VGND VGND VPWR VPWR nSEL0 sky130_fd_sc_hd__inv_2
x2 SEL1 VGND VGND VPWR VPWR nSEL1 sky130_fd_sc_hd__inv_2
x7 nSEL0 nSEL1 VGND VGND VPWR VPWR gno0 sky130_fd_sc_hd__and2_1
x10 SEL1 SEL0 VGND VGND VPWR VPWR gno3 sky130_fd_sc_hd__and2_1
x11 gno0 VGND VGND VPWR VPWR gpo0 sky130_fd_sc_hd__inv_2
x12 gno1 VGND VGND VPWR VPWR gpo1 sky130_fd_sc_hd__inv_2
x13 gno2 VGND VGND VPWR VPWR gpo2 sky130_fd_sc_hd__inv_2
x14 gno3 VGND VGND VPWR VPWR gpo3 sky130_fd_sc_hd__inv_2
x15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
x16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
x17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
x8 SEL1 SEL0 VGND VGND VPWR VPWR gno1 sky130_fd_sc_hd__and2b_1
x9 SEL0 SEL1 VGND VGND VPWR VPWR gno2 sky130_fd_sc_hd__and2b_1
x18 SEL2 VGND VGND VPWR VPWR nSEL2 sky130_fd_sc_hd__inv_2
x19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
.ends

**** begin user architecture code


* ngspice commands
* .options savecurrents
.param VCC = 1.8
.param SRCRES = 1k
.include stimuli_tb_mux8to1.cir
.control
save all
op
write tb_mux8to1.raw
set appendwrite
tran 200n 120u
write tb_mux8to1.raw
*quit 0
.endc



**** end user architecture code
.end
