* NGSPICE file created from passgate_parax.ext - technology: sky130A

.subckt passgate_parax A GN GP Z VDD VSS
X0 Z.t1 GN.t0 A.t0 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X1 A.t2 GP.t0 Z.t2 VDD.t1 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X2 Z.t0 GN.t1 A.t1 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X3 A.t3 GP.t1 Z.t3 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
R0 GN.n0 GN.t0 377.486
R1 GN.n0 GN.t1 374.202
R2 GN GN.n0 2.16602
R3 A.n0 A.t3 26.3998
R4 A.n0 A.t2 23.5483
R5 A.n1 A.t0 12.7127
R6 A.n1 A.t1 10.8578
R7 A.n2 A.n0 3.06895
R8 A.n2 A.n1 1.84731
R9 A A.n2 1.18948
R10 Z.n1 Z.t2 23.6581
R11 Z.n0 Z.t3 23.3739
R12 Z.n1 Z.t0 10.7528
R13 Z.n3 Z.t1 10.6417
R14 Z.n2 Z.n1 1.30064
R15 Z Z.n4 0.958687
R16 Z.n2 Z.n0 0.726502
R17 Z.n3 Z.n2 0.512491
R18 Z.n4 Z.n3 0.359663
R19 Z.n4 Z.n0 0.216071
R20 VSS.n6 VSS.n4 11744.7
R21 VSS.n8 VSS.n4 11744.7
R22 VSS.n8 VSS.n3 11744.7
R23 VSS.n6 VSS.n3 11744.7
R24 VSS.t1 VSS.n3 8583.05
R25 VSS.t0 VSS.n4 8583.05
R26 VSS.n7 VSS.t1 7967.33
R27 VSS.n7 VSS.t0 7967.33
R28 VSS.n5 VSS.n2 763.09
R29 VSS.n5 VSS.n0 732.236
R30 VSS.n9 VSS.n2 304.553
R31 VSS.n10 VSS.n9 266.349
R32 VSS.n3 VSS.n2 195
R33 VSS.n4 VSS.n1 195
R34 VSS.n10 VSS.n1 54.2123
R35 VSS.n1 VSS.n0 30.8711
R36 VSS.n6 VSS.n5 11.0382
R37 VSS.n7 VSS.n6 11.0382
R38 VSS.n9 VSS.n8 11.0382
R39 VSS.n8 VSS.n7 11.0382
R40 VSS.n11 VSS.n0 10.4476
R41 VSS VSS.n11 7.23036
R42 VSS.n11 VSS.n10 3.78485
R43 GP.n0 GP.t1 450.938
R44 GP.n0 GP.t0 445.666
R45 GP GP.n0 3.23793
R46 VDD.n8 VDD.n2 8629.41
R47 VDD.n8 VDD.n3 8629.41
R48 VDD.n6 VDD.n2 8629.41
R49 VDD.n6 VDD.n3 8629.41
R50 VDD.n8 VDD.t0 2459.29
R51 VDD.t1 VDD.n6 2459.29
R52 VDD.t0 VDD.n7 2298.92
R53 VDD.n7 VDD.t1 2298.92
R54 VDD.n5 VDD.n4 920.471
R55 VDD.n4 VDD.n0 914.447
R56 VDD.n5 VDD.n1 480.764
R57 VDD.n10 VDD.n1 379.2
R58 VDD.n11 VDD.n0 105.788
R59 VDD.n10 VDD.n9 63.3551
R60 VDD.n6 VDD.n5 61.6672
R61 VDD.n9 VDD.n8 61.6672
R62 VDD VDD.n11 7.60782
R63 VDD.n9 VDD.n0 6.02403
R64 VDD.n11 VDD.n10 5.18145
R65 VDD.n3 VDD.n1 2.84665
R66 VDD.n7 VDD.n3 2.84665
R67 VDD.n4 VDD.n2 2.84665
R68 VDD.n7 VDD.n2 2.84665
C0 GP A 3.81669f
C1 GN A 3.41095f
C2 GP GN 0.095282f
C3 VDD A 1.49242f
C4 GP VDD 1.13434f
C5 VDD GN 0.070087f
C6 Z A 4.51796f
C7 Z GP 0.278468f
C8 Z GN 0.415871f
C9 Z VDD 2.3841f
C10 GN VSS 3.479814f
C11 Z VSS 2.587187f
C12 GP VSS 2.214615f
C13 A VSS 4.2026f
C14 VDD VSS 9.990746f
C15 VDD.n0 VSS 0.041049f
C16 VDD.n1 VSS 0.13325f
C17 VDD.n2 VSS 0.064566f
C18 VDD.n3 VSS 0.064566f
C19 VDD.n4 VSS 0.064356f
C20 VDD.n5 VSS 0.089219f
C21 VDD.n6 VSS 0.287635f
C22 VDD.t1 VSS 0.415127f
C23 VDD.n7 VSS 0.400805f
C24 VDD.t0 VSS 0.415127f
C25 VDD.n8 VSS 0.287635f
C26 VDD.n9 VSS 0.002528f
C27 VDD.n10 VSS 0.070642f
C28 VDD.n11 VSS 0.021449f
C29 GP.t0 VSS 0.508073f
C30 GP.t1 VSS 0.522241f
C31 GP.n0 VSS 1.91856f
C32 Z.t3 VSS 0.452527f
C33 Z.n0 VSS 0.562808f
C34 Z.t2 VSS 0.464987f
C35 Z.t0 VSS 0.350399f
C36 Z.n1 VSS 2.34646f
C37 Z.n2 VSS 0.793945f
C38 Z.t1 VSS 0.343504f
C39 Z.n3 VSS 0.512912f
C40 Z.n4 VSS 0.705679f
C41 A.t3 VSS 0.768569f
C42 A.t2 VSS 0.543692f
C43 A.n0 VSS 4.21525f
C44 A.t0 VSS 0.742571f
C45 A.t1 VSS 0.426296f
C46 A.n1 VSS 4.13493f
C47 A.n2 VSS 0.675541f
C48 GN.t0 VSS 0.41457f
C49 GN.t1 VSS 0.404568f
C50 GN.n0 VSS 1.85301f
.ends

