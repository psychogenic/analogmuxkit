* NGSPICE file created from mux8to1_parax.ext - technology: sky130A

.subckt mux8to1_parax select1 select2 A1 A3 A2 A4 Z A8 select0 A7 A6 VDD A5 VSS
X0 a_5645_5909# a_5645_6085# a_5671_6037# VSS.t21 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X1 VSS.t1 select1.t0 a_5645_6085# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 x5.A select2.t0 Z.t1 VDD.t5 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X3 x4.A x3.GN1.t2 A5.t2 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X4 VSS.t49 a_5645_6461# x3.GN3 VSS.t48 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X5 x3.GP4.t3 x3.GN4.t2 VSS.t30 VSS.t29 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X6 x5.GN select2.t1 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VSS.t63 a_5645_5909# x3.GN2 VSS.t62 sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.169 ps=1.82 w=0.65 l=0.15
X8 VDD.t78 select0.t0 x1.nSEL0 VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 x5.A select2.t2 Z.t0 VDD.t2 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X10 A1.t1 x3.GP1.t4 x5.A VDD.t45 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X11 x5.A x3.GN2 A2.t2 VSS.t31 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X12 VDD.t72 VSS.t76 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X13 x4.A x5.GN Z.t7 VDD.t76 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X14 x1.nSEL0 select0.t1 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 x5.A x3.GN4.t3 A4.t1 VSS.t57 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X16 VSS.t41 VDD.t79 VSS.t40 VSS.t39 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X17 a_5671_6037# select0.t2 VSS.t43 VSS.t42 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X18 A7.t3 x3.GP3 x4.A VDD.t41 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X19 x4.A x5.GN Z.t6 VDD.t75 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X20 Z.t5 x5.GN x5.A VSS.t74 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X21 A3.t3 x3.GP3 x5.A VDD.t42 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X22 VSS.t56 select1.t1 x1.nSEL1 VSS.t55 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 x3.GP4.t1 x3.GN4.t4 VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X24 Z.t3 select2.t3 x4.A VSS.t75 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X25 VSS.t45 a_5645_7149# x3.GN4.t1 VSS.t44 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X26 VDD.t16 a_5645_6637# a_5645_6461# VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X27 x4.A x3.GN2 A6.t2 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X28 a_5645_7149# select1.t2 a_5699_7287# VSS.t64 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X29 x4.A x3.GN1.t3 A5.t1 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X30 a_5645_6637# select0.t3 VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X31 VSS.t16 x3.GN1.t4 x3.GP1.t3 VSS.t15 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 a_5699_7287# select0.t4 VSS.t61 VSS.t60 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X33 VSS.t68 VDD.t80 VSS.t67 VSS.t66 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X34 x5.A x3.GN3 A3.t1 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X35 A8.t3 x3.GP4.t4 x4.A VDD.t22 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X36 A1.t0 x3.GP1.t5 x5.A VDD.t45 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X37 a_5645_6461# a_5645_6637# a_5671_6589# VSS.t17 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0504 ps=0.66 w=0.42 l=0.15
X38 x5.A x3.GN4.t5 A4.t0 VSS.t57 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X39 VSS.t12 x3.GN3 x3.GP3 VSS.t11 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X40 x3.GP1.t2 x3.GN1.t5 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X41 VSS.t24 select0.t5 a_5645_6637# VSS.t23 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X42 Z.t4 x5.GN x5.A VSS.t73 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X43 VDD.t58 select1.t3 x1.nSEL1 VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X44 VDD.t56 select1.t4 a_5645_7149# VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X45 A5.t3 x3.GP1.t6 x4.A VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X46 VDD.t69 VSS.t77 VDD.t68 VDD.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X47 Z.t2 select2.t4 x4.A VSS.t65 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X48 VDD.t38 a_5645_5493# x3.GN1.t0 VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X49 a_5645_7149# select0.t6 VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X50 VDD.t74 x3.GN1.t6 x3.GP1.t1 VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X51 x4.A x3.GN3 A7.t1 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X52 x4.A x3.GN2 A6.t1 VSS.t36 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X53 A4.t3 x3.GP4.t5 x5.A VDD.t10 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X54 VSS.t70 select2.t5 x5.GN VSS.t69 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 a_5645_5493# x1.nSEL0 a_5699_5631# VSS.t54 sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X56 x1.nSEL1 select1.t5 VSS.t38 VSS.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X57 x5.A x3.GN1.t7 A1.t3 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X58 VDD.t14 x3.GN3 x3.GP3 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X59 x3.GP1.t0 x3.GN1.t8 VDD.t26 VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X60 a_5645_5909# select0.t7 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X61 x5.A x3.GN3 A3.t0 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X62 A2.t3 x3.GP2.t4 x5.A VDD.t17 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X63 x5.A x3.GN1.t9 A1.t2 VSS.t26 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X64 A3.t2 x3.GP3 x5.A VDD.t42 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X65 VDD.t66 VSS.t78 VDD.t65 VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X66 a_5699_5631# x1.nSEL1 VSS.t53 VSS.t52 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X67 VSS.t20 VDD.t81 VSS.t19 VSS.t18 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X68 x4.A x3.GN4.t6 A8.t1 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X69 VDD.t40 a_5645_6461# x3.GN3 VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X70 VSS.t35 x3.GN2 x3.GP2.t3 VSS.t34 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X71 A6.t0 x3.GP2.t5 x4.A VDD.t7 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X72 A5.t0 x3.GP1.t7 x4.A VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X73 VDD.t47 x1.nSEL0 a_5645_5493# VDD.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X74 x3.GP2.t2 x3.GN2 VSS.t33 VSS.t32 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X75 VSS.t14 x3.GN4.t7 x3.GP4.t2 VSS.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X76 VDD.t60 a_5645_5909# x3.GN2 VDD.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.26 ps=2.52 w=1 l=0.15
X77 x3.GP3 x3.GN3 VSS.t9 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X78 A7.t2 x3.GP3 x4.A VDD.t41 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X79 x1.nSEL1 select1.t6 VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X80 VDD.t1 select2.t6 x5.GN VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X81 a_5671_6589# select1.t7 VSS.t72 VSS.t71 sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1013 ps=0.99 w=0.42 l=0.15
X82 x4.A x3.GN3 A7.t0 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X83 A8.t2 x3.GP4.t6 x4.A VDD.t22 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X84 A4.t2 x3.GP4.t7 x5.A VDD.t10 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X85 a_5645_5493# x1.nSEL1 VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.16655 ps=1.39 w=0.42 l=0.15
X86 VSS.t47 a_5645_5493# x3.GN1.t1 VSS.t46 sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X87 VSS.t4 VDD.t82 VSS.t3 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X88 x5.A x3.GN2 A2.t1 VSS.t31 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X89 VDD.t32 x3.GN2 x3.GP2.t1 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X90 A2.t0 x3.GP2.t6 x5.A VDD.t17 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
X91 VDD.t36 a_5645_7149# x3.GN4.t0 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.475 ps=2.95 w=1 l=0.15
X92 x5.GN select2.t7 VSS.t28 VSS.t27 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X93 VSS.t59 select0.t8 x1.nSEL0 VSS.t58 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X94 x3.GP2.t0 x3.GN2 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X95 VDD.t34 x3.GN4.t8 x3.GP4.t0 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X96 x4.A x3.GN4.t9 A8.t0 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=0.35
X97 VDD.t21 a_5645_6085# a_5645_5909# VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.0609 ps=0.71 w=0.42 l=0.15
X98 x3.GP3 x3.GN3 VDD.t12 VDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X99 VDD.t63 VSS.t79 VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X100 a_5645_6085# select1.t8 VDD.t52 VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0714 ps=0.76 w=0.42 l=0.15
X101 x1.nSEL0 select0.t9 VSS.t51 VSS.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X102 a_5645_6461# select1.t9 VDD.t50 VDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.2279 ps=1.74 w=0.42 l=0.15
X103 A6.t3 x3.GP2.t7 x4.A VDD.t7 sky130_fd_pr__pfet_01v8_lvt ad=2.9 pd=20.58 as=2.9 ps=20.58 w=10 l=0.35
R0 VSS.n163 VSS.n162 587674
R1 VSS.n219 VSS.n218 153375
R2 VSS.n119 VSS.n112 117542
R3 VSS.n177 VSS.n176 71206.2
R4 VSS.n176 VSS.n175 64736.2
R5 VSS.n164 VSS.n9 16580.8
R6 VSS.n168 VSS.n108 11744.7
R7 VSS.n174 VSS.n108 11744.7
R8 VSS.n168 VSS.n109 11744.7
R9 VSS.n174 VSS.n109 11744.7
R10 VSS.n116 VSS.n106 11744.7
R11 VSS.n178 VSS.n106 11744.7
R12 VSS.n116 VSS.n107 11744.7
R13 VSS.n178 VSS.n107 11744.7
R14 VSS.n267 VSS.n22 11744.7
R15 VSS.n263 VSS.n22 11744.7
R16 VSS.n267 VSS.n23 11744.7
R17 VSS.n263 VSS.n23 11744.7
R18 VSS.n281 VSS.n10 11744.7
R19 VSS.n277 VSS.n10 11744.7
R20 VSS.n281 VSS.n11 11744.7
R21 VSS.n277 VSS.n11 11744.7
R22 VSS.n274 VSS.n16 11744.7
R23 VSS.n270 VSS.n16 11744.7
R24 VSS.n274 VSS.n17 11744.7
R25 VSS.n270 VSS.n17 11744.7
R26 VSS.n256 VSS.n28 11744.7
R27 VSS.n256 VSS.n29 11744.7
R28 VSS.n260 VSS.n29 11744.7
R29 VSS.n260 VSS.n28 11744.7
R30 VSS.n131 VSS.n130 11744.7
R31 VSS.n127 VSS.n126 11744.7
R32 VSS.n130 VSS.n127 11744.7
R33 VSS.n160 VSS.n120 11744.7
R34 VSS.n156 VSS.n121 11744.7
R35 VSS.n160 VSS.n121 11744.7
R36 VSS.n144 VSS.n143 11744.7
R37 VSS.n140 VSS.n139 11744.7
R38 VSS.n143 VSS.n140 11744.7
R39 VSS.n284 VSS.n4 11744.7
R40 VSS.n284 VSS.n5 11744.7
R41 VSS.n7 VSS.n4 11744.7
R42 VSS.n163 VSS.n112 10428.2
R43 VSS.n164 VSS.n117 7573.12
R44 VSS.n117 VSS.t73 7065.1
R45 VSS.n177 VSS.t74 7065.1
R46 VSS.t73 VSS.n113 6710.74
R47 VSS.n113 VSS.t74 6710.74
R48 VSS.n167 VSS.n165 6647.5
R49 VSS.n276 VSS.n275 6049.9
R50 VSS.n167 VSS.t75 6006.85
R51 VSS.n175 VSS.t65 6006.85
R52 VSS.n262 VSS.n261 6004.3
R53 VSS.n283 VSS.n282 5972.7
R54 VSS.n269 VSS.n268 5963.12
R55 VSS.t75 VSS.n166 5705.56
R56 VSS.n166 VSS.t65 5705.56
R57 VSS.n165 VSS.n112 4796.58
R58 VSS.n164 VSS.n163 3666.67
R59 VSS.n118 VSS.n9 3385.09
R60 VSS.n15 VSS.n9 3361.58
R61 VSS.n27 VSS.n21 3305.56
R62 VSS.n161 VSS.n119 3279.94
R63 VSS.n21 VSS.n15 3275.35
R64 VSS.n68 VSS.n27 2366.85
R65 VSS.n176 VSS.n33 2235.82
R66 VSS.n162 VSS.n161 1652.78
R67 VSS.n162 VSS.n118 1652.78
R68 VSS.t44 VSS.n57 1550.96
R69 VSS VSS.t23 1289.66
R70 VSS.n82 VSS.n69 1198.25
R71 VSS.n222 VSS.n220 1198.25
R72 VSS.n231 VSS.n57 1194.5
R73 VSS.n252 VSS.n251 1171.32
R74 VSS.n254 VSS.n33 1006.48
R75 VSS VSS.n57 918.774
R76 VSS.t46 VSS 918.774
R77 VSS.t60 VSS.t44 910.346
R78 VSS.t71 VSS.t48 826.054
R79 VSS.t42 VSS.t62 826.054
R80 VSS.t0 VSS.t55 792.337
R81 VSS.n273 VSS.n272 767.294
R82 VSS.n259 VSS.n258 767.294
R83 VSS.n158 VSS.n157 767.294
R84 VSS.n6 VSS.n3 767.294
R85 VSS.n266 VSS.n265 763.106
R86 VSS.n280 VSS.n279 763.106
R87 VSS.n128 VSS.n124 763.106
R88 VSS.n141 VSS.n137 763.106
R89 VSS.n169 VSS.n111 763.09
R90 VSS.n115 VSS.n105 763.09
R91 VSS.n111 VSS.n110 732.236
R92 VSS.n266 VSS.n24 732.236
R93 VSS.n280 VSS.n12 732.236
R94 VSS.n273 VSS.n18 732.236
R95 VSS.n259 VSS.n30 732.236
R96 VSS.n180 VSS.n105 732.236
R97 VSS.n133 VSS.n124 732.236
R98 VSS.n157 VSS.n154 732.236
R99 VSS.n146 VSS.n137 732.236
R100 VSS.n6 VSS.n1 732.236
R101 VSS.n219 VSS.n33 709.912
R102 VSS.t69 VSS.t27 708.047
R103 VSS.t55 VSS.t37 708.047
R104 VSS.t58 VSS.t50 708.047
R105 VSS.t54 VSS.t52 708.047
R106 VSS.t39 VSS.n252 606.351
R107 VSS.t64 VSS 564.751
R108 VSS.t27 VSS 564.751
R109 VSS.t50 VSS 564.751
R110 VSS VSS.t54 564.751
R111 VSS VSS.n219 564.751
R112 VSS.n218 VSS.t64 522.606
R113 VSS.t52 VSS.t18 522.606
R114 VSS.t21 VSS 480.461
R115 VSS VSS.t2 408.628
R116 VSS.t18 VSS.t46 387.74
R117 VSS VSS.n253 384.901
R118 VSS.n69 VSS.t34 374.356
R119 VSS.n220 VSS.t17 337.166
R120 VSS.n255 VSS.n254 332.642
R121 VSS.t13 VSS 329.539
R122 VSS.t11 VSS 329.539
R123 VSS VSS.t15 329.539
R124 VSS.n272 VSS.n271 325.502
R125 VSS.n258 VSS.n257 325.502
R126 VSS.n159 VSS.n158 325.502
R127 VSS.n285 VSS.n3 325.502
R128 VSS.n220 VSS.t71 320.307
R129 VSS.n170 VSS.n169 304.553
R130 VSS.n115 VSS.n114 304.553
R131 VSS.n265 VSS.n264 304.204
R132 VSS.n279 VSS.n278 304.204
R133 VSS.n129 VSS.n128 304.204
R134 VSS.n142 VSS.n141 304.204
R135 VSS.t17 VSS 295.019
R136 VSS.n172 VSS.n170 266.349
R137 VSS.n114 VSS.n104 266.349
R138 VSS VSS.t0 261.303
R139 VSS.t66 VSS 244.445
R140 VSS.n264 VSS.n26 242.448
R141 VSS.n278 VSS.n14 242.448
R142 VSS.n271 VSS.n20 242.448
R143 VSS.n257 VSS.n32 242.448
R144 VSS.n129 VSS.n123 242.448
R145 VSS.n159 VSS.n122 242.448
R146 VSS.n142 VSS.n136 242.448
R147 VSS.n286 VSS.n285 242.448
R148 VSS.n238 VSS.t1 240.575
R149 VSS.n216 VSS.t24 237.327
R150 VSS.t29 VSS.t13 221.451
R151 VSS.t8 VSS.t11 221.451
R152 VSS.t34 VSS.t32 221.451
R153 VSS.t15 VSS.t5 221.451
R154 VSS.n195 VSS.t79 218.308
R155 VSS.n61 VSS.t78 218.308
R156 VSS.n42 VSS.t77 218.308
R157 VSS.n225 VSS.t76 218.308
R158 VSS.n192 VSS.t40 214.456
R159 VSS.n194 VSS.t41 214.456
R160 VSS.n205 VSS.t3 214.456
R161 VSS.n62 VSS.t4 214.456
R162 VSS.n37 VSS.t19 214.456
R163 VSS.n41 VSS.t20 214.456
R164 VSS.n230 VSS.t67 214.456
R165 VSS.n224 VSS.t68 214.456
R166 VSS.n210 VSS.n209 204.457
R167 VSS.n50 VSS.n49 200.231
R168 VSS.n55 VSS.n54 200.231
R169 VSS.n44 VSS.n39 200.105
R170 VSS.n69 VSS 197.724
R171 VSS.n252 VSS 197.724
R172 VSS.n272 VSS.n17 195
R173 VSS.n17 VSS.t10 195
R174 VSS.n19 VSS.n16 195
R175 VSS.n16 VSS.t10 195
R176 VSS.n279 VSS.n11 195
R177 VSS.n11 VSS.t57 195
R178 VSS.n13 VSS.n10 195
R179 VSS.n10 VSS.t57 195
R180 VSS.n265 VSS.n23 195
R181 VSS.n23 VSS.t31 195
R182 VSS.n25 VSS.n22 195
R183 VSS.n22 VSS.t31 195
R184 VSS.n31 VSS.n28 195
R185 VSS.n253 VSS.n28 195
R186 VSS.n258 VSS.n29 195
R187 VSS.n29 VSS.t26 195
R188 VSS.n179 VSS.n178 195
R189 VSS.n178 VSS.n177 195
R190 VSS.n116 VSS.n115 195
R191 VSS.n117 VSS.n116 195
R192 VSS.n174 VSS.n173 195
R193 VSS.n175 VSS.n174 195
R194 VSS.n169 VSS.n168 195
R195 VSS.n168 VSS.n167 195
R196 VSS.n128 VSS.n127 195
R197 VSS.n127 VSS.t25 195
R198 VSS.n132 VSS.n131 195
R199 VSS.n158 VSS.n121 195
R200 VSS.n121 VSS.t7 195
R201 VSS.n153 VSS.n120 195
R202 VSS.n141 VSS.n140 195
R203 VSS.n140 VSS.t36 195
R204 VSS.n145 VSS.n144 195
R205 VSS.n4 VSS.n2 195
R206 VSS.t22 VSS.n4 195
R207 VSS.n5 VSS.n3 195
R208 VSS.n8 VSS.n5 188.989
R209 VSS.n144 VSS.n138 188.988
R210 VSS.n155 VSS.n120 188.986
R211 VSS.n131 VSS.n125 188.984
R212 VSS.n218 VSS.t60 185.441
R213 VSS.n261 VSS.t26 183.936
R214 VSS VSS.t42 177.012
R215 VSS VSS.t8 176.633
R216 VSS.t32 VSS 176.633
R217 VSS.t5 VSS 176.633
R218 VSS.n254 VSS 176.633
R219 VSS.n126 VSS.n125 173.373
R220 VSS.n156 VSS.n155 173.304
R221 VSS.n139 VSS.n138 173.167
R222 VSS.n8 VSS.n7 173.097
R223 VSS.n90 VSS.t14 162.471
R224 VSS.n85 VSS.t12 162.471
R225 VSS.n81 VSS.t35 162.471
R226 VSS.n76 VSS.t16 162.471
R227 VSS.n239 VSS.t56 162.471
R228 VSS.n50 VSS.t59 160.046
R229 VSS.n55 VSS.t70 160.046
R230 VSS.n64 VSS.t30 160.017
R231 VSS.n83 VSS.t9 160.017
R232 VSS.n71 VSS.t33 160.017
R233 VSS.n74 VSS.t6 160.017
R234 VSS.n246 VSS.t51 160.017
R235 VSS.n241 VSS.t38 160.017
R236 VSS.n238 VSS.t28 158.534
R237 VSS.n275 VSS.t10 155.954
R238 VSS.n282 VSS.t57 155.954
R239 VSS.n268 VSS.t31 155.831
R240 VSS.n255 VSS.t26 139.648
R241 VSS.n130 VSS.n119 118.54
R242 VSS.n161 VSS.n160 111.895
R243 VSS.n143 VSS.n118 111.808
R244 VSS.n276 VSS.n15 99.881
R245 VSS.n269 VSS.n21 93.748
R246 VSS.n262 VSS.n27 93.6734
R247 VSS.n68 VSS.t29 89.635
R248 VSS.n9 VSS.t22 89.4314
R249 VSS VSS.n68 86.9987
R250 VSS.t37 VSS.t21 84.2917
R251 VSS.n165 VSS.n164 79.0175
R252 VSS.n39 VSS.t53 72.8576
R253 VSS.n209 VSS.t61 72.8576
R254 VSS.n283 VSS.n9 72.6343
R255 VSS.n161 VSS.t7 66.9242
R256 VSS.t36 VSS.n118 66.8669
R257 VSS.n21 VSS.t10 62.2068
R258 VSS.n27 VSS.t31 62.1573
R259 VSS.t25 VSS.n119 60.352
R260 VSS.n49 VSS.t43 58.5719
R261 VSS.n54 VSS.t72 58.5719
R262 VSS.n15 VSS.t57 56.0738
R263 VSS.n173 VSS.n172 54.2123
R264 VSS.n179 VSS.n104 54.2123
R265 VSS.t48 VSS.t69 50.5752
R266 VSS.t62 VSS.t58 50.5752
R267 VSS.n208 VSS 43.9579
R268 VSS.n256 VSS.n255 42.2329
R269 VSS.n211 VSS.n208 34.6358
R270 VSS.n215 VSS.n58 34.6358
R271 VSS.n173 VSS.n110 30.8711
R272 VSS.n25 VSS.n24 30.8711
R273 VSS.n13 VSS.n12 30.8711
R274 VSS.n19 VSS.n18 30.8711
R275 VSS.n31 VSS.n30 30.8711
R276 VSS.n180 VSS.n179 30.8711
R277 VSS.n133 VSS.n132 30.8711
R278 VSS.n154 VSS.n153 30.8711
R279 VSS.n146 VSS.n145 30.8711
R280 VSS.n2 VSS.n1 30.8711
R281 VSS.n251 VSS.n34 26.9246
R282 VSS.n231 VSS.n215 25.6926
R283 VSS.n49 VSS.t63 25.4291
R284 VSS.n54 VSS.t49 25.4291
R285 VSS.n90 VSS.n89 25.224
R286 VSS.n89 VSS.n64 25.224
R287 VSS.n85 VSS.n84 25.224
R288 VSS.n84 VSS.n83 25.224
R289 VSS.n81 VSS.n80 25.224
R290 VSS.n80 VSS.n71 25.224
R291 VSS.n76 VSS.n75 25.224
R292 VSS.n75 VSS.n74 25.224
R293 VSS.n246 VSS.n245 25.224
R294 VSS.n240 VSS.n239 25.224
R295 VSS.n241 VSS.n240 25.224
R296 VSS.n238 VSS.n237 24.0946
R297 VSS.n253 VSS.t39 23.7273
R298 VSS.n39 VSS.t47 22.3257
R299 VSS.n209 VSS.t45 22.3257
R300 VSS.n245 VSS.n50 21.4593
R301 VSS.n237 VSS.n55 21.4593
R302 VSS.n85 VSS.n64 20.3299
R303 VSS.n76 VSS.n71 20.3299
R304 VSS.n91 VSS.n90 19.2926
R305 VSS.n246 VSS.n48 17.7867
R306 VSS.n82 VSS.n81 17.3181
R307 VSS.t23 VSS.t66 16.8587
R308 VSS.n83 VSS.n82 15.8123
R309 VSS.n74 VSS.n34 15.8123
R310 VSS.n284 VSS.n283 15.1478
R311 VSS.n191 VSS.n34 14.775
R312 VSS.n223 VSS.n222 14.775
R313 VSS.n239 VSS.n238 13.5534
R314 VSS.n207 VSS.n206 11.2844
R315 VSS.n271 VSS.n270 11.0382
R316 VSS.n270 VSS.n269 11.0382
R317 VSS.n274 VSS.n273 11.0382
R318 VSS.n275 VSS.n274 11.0382
R319 VSS.n278 VSS.n277 11.0382
R320 VSS.n277 VSS.n276 11.0382
R321 VSS.n281 VSS.n280 11.0382
R322 VSS.n282 VSS.n281 11.0382
R323 VSS.n264 VSS.n263 11.0382
R324 VSS.n263 VSS.n262 11.0382
R325 VSS.n267 VSS.n266 11.0382
R326 VSS.n268 VSS.n267 11.0382
R327 VSS.n260 VSS.n259 11.0382
R328 VSS.n261 VSS.n260 11.0382
R329 VSS.n257 VSS.n256 11.0382
R330 VSS.n114 VSS.n107 11.0382
R331 VSS.n113 VSS.n107 11.0382
R332 VSS.n106 VSS.n105 11.0382
R333 VSS.n113 VSS.n106 11.0382
R334 VSS.n170 VSS.n109 11.0382
R335 VSS.n166 VSS.n109 11.0382
R336 VSS.n111 VSS.n108 11.0382
R337 VSS.n166 VSS.n108 11.0382
R338 VSS.n130 VSS.n129 11.0382
R339 VSS.n126 VSS.n124 11.0382
R340 VSS.n160 VSS.n159 11.0382
R341 VSS.n157 VSS.n156 11.0382
R342 VSS.n143 VSS.n142 11.0382
R343 VSS.n139 VSS.n137 11.0382
R344 VSS.n7 VSS.n6 11.0382
R345 VSS.n285 VSS.n284 11.0382
R346 VSS.n26 VSS.n25 10.9181
R347 VSS.n14 VSS.n13 10.9181
R348 VSS.n20 VSS.n19 10.9181
R349 VSS.n32 VSS.n31 10.9181
R350 VSS.n132 VSS.n123 10.9181
R351 VSS.n153 VSS.n122 10.9181
R352 VSS.n145 VSS.n136 10.9181
R353 VSS.n286 VSS.n2 10.9181
R354 VSS.n171 VSS.n110 10.4476
R355 VSS.n95 VSS.n24 10.4476
R356 VSS.n99 VSS.n12 10.4476
R357 VSS.n97 VSS.n18 10.4476
R358 VSS.n93 VSS.n30 10.4476
R359 VSS.n181 VSS.n180 10.4476
R360 VSS.n134 VSS.n133 10.4476
R361 VSS.n154 VSS.n152 10.4476
R362 VSS.n147 VSS.n146 10.4476
R363 VSS.n287 VSS.n1 10.4476
R364 VSS.n241 VSS.n50 10.1652
R365 VSS.n194 VSS.n189 9.70901
R366 VSS.n206 VSS.n205 9.70901
R367 VSS.n41 VSS.n40 9.70901
R368 VSS.n210 VSS.n58 9.41227
R369 VSS.n251 VSS.n250 9.3005
R370 VSS.n74 VSS.n73 9.3005
R371 VSS.n78 VSS.n71 9.3005
R372 VSS.n82 VSS.n67 9.3005
R373 VSS.n83 VSS.n66 9.3005
R374 VSS.n87 VSS.n64 9.3005
R375 VSS.n92 VSS.n91 9.3005
R376 VSS.n203 VSS.n202 9.3005
R377 VSS.n204 VSS.n60 9.3005
R378 VSS.n90 VSS.n63 9.3005
R379 VSS.n89 VSS.n88 9.3005
R380 VSS.n86 VSS.n85 9.3005
R381 VSS.n84 VSS.n65 9.3005
R382 VSS.n81 VSS.n70 9.3005
R383 VSS.n80 VSS.n79 9.3005
R384 VSS.n77 VSS.n76 9.3005
R385 VSS.n75 VSS.n72 9.3005
R386 VSS.n197 VSS.n196 9.3005
R387 VSS.n193 VSS.n188 9.3005
R388 VSS.n191 VSS.n190 9.3005
R389 VSS.n36 VSS.n34 9.3005
R390 VSS.n232 VSS.n231 9.3005
R391 VSS.n229 VSS.n228 9.3005
R392 VSS.n56 VSS.n55 9.3005
R393 VSS.n238 VSS.n53 9.3005
R394 VSS.n243 VSS.n50 9.3005
R395 VSS.n43 VSS.n38 9.3005
R396 VSS.n46 VSS.n45 9.3005
R397 VSS.n48 VSS.n47 9.3005
R398 VSS.n247 VSS.n246 9.3005
R399 VSS.n245 VSS.n244 9.3005
R400 VSS.n242 VSS.n241 9.3005
R401 VSS.n240 VSS.n51 9.3005
R402 VSS.n239 VSS.n52 9.3005
R403 VSS.n237 VSS.n236 9.3005
R404 VSS.n223 VSS.n217 9.3005
R405 VSS.n227 VSS.n226 9.3005
R406 VSS.n215 VSS.n214 9.3005
R407 VSS.n213 VSS.n58 9.3005
R408 VSS.n212 VSS.n211 9.3005
R409 VSS.n208 VSS.n59 9.3005
R410 VSS.n222 VSS.n221 9.3005
R411 VSS.n101 VSS.n100 8.45078
R412 VSS.n150 VSS.n135 8.45078
R413 VSS.n184 VSS.n94 8.30267
R414 VSS.n288 VSS.n0 8.30267
R415 VSS.n102 VSS.n96 7.97888
R416 VSS.n149 VSS.n148 7.97888
R417 VSS.n101 VSS.n98 7.97601
R418 VSS.n151 VSS.n150 7.97601
R419 VSS.n171 VSS.n103 7.16724
R420 VSS.n96 VSS.n95 7.16724
R421 VSS.n100 VSS.n99 7.16724
R422 VSS.n98 VSS.n97 7.16724
R423 VSS.n94 VSS.n93 7.16724
R424 VSS.n182 VSS.n181 7.16724
R425 VSS.n135 VSS.n134 7.16724
R426 VSS.n152 VSS.n151 7.16724
R427 VSS.n148 VSS.n147 7.16724
R428 VSS.n288 VSS.n287 7.16724
R429 VSS.n222 VSS.n55 7.15344
R430 VSS.n249 VSS.n248 6.50373
R431 VSS.n211 VSS.n210 6.4005
R432 VSS.n196 VSS.n193 6.26433
R433 VSS.n204 VSS.n203 6.26433
R434 VSS.n193 VSS.n192 5.85582
R435 VSS.n205 VSS.n204 5.85582
R436 VSS.n45 VSS.n37 5.85582
R437 VSS.n230 VSS.n229 5.85582
R438 VSS.n226 VSS.n216 5.85582
R439 VSS.n249 VSS.n36 4.788
R440 VSS.n95 VSS.n26 4.73093
R441 VSS.n99 VSS.n14 4.73093
R442 VSS.n97 VSS.n20 4.73093
R443 VSS.n93 VSS.n32 4.73093
R444 VSS.n134 VSS.n123 4.73093
R445 VSS.n152 VSS.n122 4.73093
R446 VSS.n147 VSS.n136 4.73093
R447 VSS.n287 VSS.n286 4.73093
R448 VSS.n250 VSS.n249 4.50726
R449 VSS.n186 VSS 4.01425
R450 VSS.n185 VSS 4.01425
R451 VSS.n172 VSS.n171 3.78485
R452 VSS.n181 VSS.n104 3.78485
R453 VSS.n44 VSS.n43 3.40476
R454 VSS.n196 VSS.n195 3.13241
R455 VSS.n203 VSS.n61 3.13241
R456 VSS.n43 VSS.n42 3.13241
R457 VSS.n226 VSS.n225 3.13241
R458 VSS.n234 VSS.n233 2.88636
R459 VSS.t25 VSS.n125 2.87953
R460 VSS.n155 VSS.t7 2.87839
R461 VSS.t36 VSS.n138 2.87611
R462 VSS.t22 VSS.n8 2.87497
R463 VSS.n45 VSS.n44 2.86007
R464 VSS.n195 VSS.n194 2.7239
R465 VSS.n62 VSS.n61 2.7239
R466 VSS.n42 VSS.n41 2.7239
R467 VSS.n225 VSS.n224 2.7239
R468 VSS.n183 VSS.n103 2.03666
R469 VSS.n183 VSS.n182 1.77451
R470 VSS.n201 VSS.n200 1.753
R471 VSS.n199 VSS.n198 1.753
R472 VSS VSS.n187 1.48125
R473 VSS.n184 VSS.n183 1.44312
R474 VSS.n235 VSS.n234 1.21169
R475 VSS.n187 VSS.n186 1.11894
R476 VSS.n200 VSS 0.95037
R477 VSS.n200 VSS.n199 0.761313
R478 VSS.n234 VSS 0.531208
R479 VSS.n102 VSS.n101 0.467019
R480 VSS.n150 VSS.n149 0.467019
R481 VSS.n192 VSS.n191 0.409011
R482 VSS.n91 VSS.n62 0.409011
R483 VSS.n48 VSS.n37 0.409011
R484 VSS.n231 VSS.n230 0.409011
R485 VSS.n229 VSS.n216 0.409011
R486 VSS.n224 VSS.n223 0.409011
R487 VSS.n186 VSS.n0 0.198729
R488 VSS.n185 VSS.n184 0.194976
R489 VSS.n250 VSS.n35 0.1255
R490 VSS.n206 VSS.n60 0.120292
R491 VSS.n202 VSS.n60 0.120292
R492 VSS.n88 VSS.n63 0.120292
R493 VSS.n88 VSS.n87 0.120292
R494 VSS.n86 VSS.n65 0.120292
R495 VSS.n66 VSS.n65 0.120292
R496 VSS.n79 VSS.n70 0.120292
R497 VSS.n79 VSS.n78 0.120292
R498 VSS.n77 VSS.n72 0.120292
R499 VSS.n73 VSS.n72 0.120292
R500 VSS.n190 VSS.n188 0.120292
R501 VSS.n197 VSS.n189 0.120292
R502 VSS.n212 VSS.n59 0.120292
R503 VSS.n213 VSS.n212 0.120292
R504 VSS.n214 VSS.n213 0.120292
R505 VSS.n227 VSS.n217 0.120292
R506 VSS.n52 VSS.n51 0.120292
R507 VSS.n242 VSS.n51 0.120292
R508 VSS.n244 VSS.n243 0.120292
R509 VSS.n47 VSS.n46 0.120292
R510 VSS.n46 VSS.n38 0.120292
R511 VSS.n40 VSS.n38 0.120292
R512 VSS VSS.n227 0.0981562
R513 VSS VSS.n207 0.09425
R514 VSS.n199 VSS 0.0881354
R515 VSS.n184 VSS.n102 0.0766574
R516 VSS.n149 VSS.n0 0.0766574
R517 VSS.n198 VSS.n197 0.0721146
R518 VSS.n236 VSS.n235 0.0708125
R519 VSS.n96 VSS 0.064875
R520 VSS.n98 VSS 0.064875
R521 VSS.n94 VSS 0.064875
R522 VSS.n151 VSS 0.064875
R523 VSS.n148 VSS 0.064875
R524 VSS VSS.n288 0.064875
R525 VSS.n100 VSS 0.063625
R526 VSS.n135 VSS 0.063625
R527 VSS.n202 VSS.n201 0.0616979
R528 VSS.n103 VSS 0.061125
R529 VSS.n182 VSS 0.061125
R530 VSS.n63 VSS 0.0603958
R531 VSS VSS.n86 0.0603958
R532 VSS.n67 VSS 0.0603958
R533 VSS.n70 VSS 0.0603958
R534 VSS VSS.n77 0.0603958
R535 VSS VSS.n36 0.0603958
R536 VSS.n190 VSS 0.0603958
R537 VSS.n214 VSS 0.0603958
R538 VSS.n228 VSS 0.0603958
R539 VSS.n221 VSS 0.0603958
R540 VSS VSS.n56 0.0603958
R541 VSS.n236 VSS 0.0603958
R542 VSS VSS.n53 0.0603958
R543 VSS VSS.n52 0.0603958
R544 VSS.n243 VSS 0.0603958
R545 VSS.n244 VSS 0.0603958
R546 VSS.n47 VSS 0.0603958
R547 VSS.n201 VSS.n92 0.0590938
R548 VSS.n248 VSS 0.0590938
R549 VSS.n235 VSS.n56 0.0499792
R550 VSS.n198 VSS.n188 0.0486771
R551 VSS.n233 VSS 0.0460729
R552 VSS.n187 VSS.n185 0.040297
R553 VSS.n232 VSS 0.0343542
R554 VSS VSS.n67 0.0330521
R555 VSS.n221 VSS 0.0330521
R556 VSS VSS.n35 0.03175
R557 VSS.n92 VSS 0.0226354
R558 VSS.n87 VSS 0.0226354
R559 VSS VSS.n66 0.0226354
R560 VSS.n78 VSS 0.0226354
R561 VSS.n73 VSS 0.0226354
R562 VSS.n189 VSS 0.0226354
R563 VSS.n228 VSS 0.0226354
R564 VSS VSS.n217 0.0226354
R565 VSS.n53 VSS 0.0226354
R566 VSS VSS.n242 0.0226354
R567 VSS.n247 VSS 0.0226354
R568 VSS.n40 VSS 0.0226354
R569 VSS.n233 VSS.n232 0.0148229
R570 VSS.n207 VSS.n59 0.00440625
R571 VSS.n36 VSS.n35 0.00180208
R572 VSS.n248 VSS.n247 0.00180208
R573 select1.n10 select1.t8 327.99
R574 select1.n3 select1.t7 293.969
R575 select1.n6 select1.t4 256.07
R576 select1.n1 select1.t6 212.081
R577 select1.n0 select1.t3 212.081
R578 select1.n10 select1.t0 199.457
R579 select1.n2 select1.n1 182.929
R580 select1 select1.n3 154.065
R581 select1.n11 select1.n10 152
R582 select1.n7 select1.n6 152
R583 select1.n6 select1.t2 150.03
R584 select1.n1 select1.t5 139.78
R585 select1.n0 select1.t1 139.78
R586 select1.n3 select1.t9 138.338
R587 select1.n1 select1.n0 61.346
R588 select1.n5 select1 22.1096
R589 select1.n14 select1.n13 14.6836
R590 select1.n13 select1.n12 14.6704
R591 select1.n12 select1 13.8672
R592 select1.n4 select1 13.8328
R593 select1.n11 select1 12.1605
R594 select1.n14 select1.n2 10.6811
R595 select1.n7 select1.n5 10.4374
R596 select1.n9 select1.n8 8.15359
R597 select1.n2 select1 6.1445
R598 select1.n4 select1 5.16179
R599 select1.n9 select1.n4 4.65206
R600 select1.n8 select1 3.93896
R601 select1 select1.n11 2.34717
R602 select1.n5 select1 2.16665
R603 select1.n8 select1.n7 1.57588
R604 select1.n13 select1.n9 0.79438
R605 select1.n12 select1 0.6405
R606 select1 select1.n14 0.248606
R607 select2.n5 select2.t0 450.938
R608 select2.n5 select2.t2 445.666
R609 select2.n0 select2.t3 377.486
R610 select2.n0 select2.t4 374.202
R611 select2.n2 select2.t1 212.081
R612 select2.n1 select2.t6 212.081
R613 select2.n3 select2.n2 183.441
R614 select2.n2 select2.t7 139.78
R615 select2.n1 select2.t5 139.78
R616 select2.n2 select2.n1 61.346
R617 select2.n8 select2.n7 12.4093
R618 select2 select2.n3 11.4331
R619 select2.n7 select2.n6 9.10647
R620 select2.n7 select2.n4 8.98648
R621 select2.n3 select2 5.6325
R622 select2.n4 select2 5.02323
R623 select2.n6 select2.n5 3.1748
R624 select2.n8 select2.n0 2.10165
R625 select2.n4 select2 0.941788
R626 select2 select2.n8 0.064875
R627 select2.n6 select2 0.063625
R628 Z.n1 Z.t0 23.6581
R629 Z.n7 Z.t7 23.6581
R630 Z.n0 Z.t1 23.3739
R631 Z.n6 Z.t6 23.3739
R632 Z.n1 Z.t5 10.7528
R633 Z.n7 Z.t2 10.7528
R634 Z.n3 Z.t4 10.6417
R635 Z.n9 Z.t3 10.6417
R636 Z.n2 Z.n1 1.30064
R637 Z.n8 Z.n7 1.30064
R638 Z.n11 Z.n10 1.04212
R639 Z Z.n5 0.919875
R640 Z.n5 Z.n4 0.859481
R641 Z.n11 Z 0.754624
R642 Z.n2 Z.n0 0.726502
R643 Z.n8 Z.n6 0.726502
R644 Z.n3 Z.n2 0.512491
R645 Z.n9 Z.n8 0.512491
R646 Z.n4 Z.n3 0.359663
R647 Z.n10 Z.n9 0.359663
R648 Z.n4 Z.n0 0.216071
R649 Z.n10 Z.n6 0.216071
R650 Z Z.n11 0.0100278
R651 Z.n5 Z 0.001125
R652 VDD.n190 VDD.n188 8629.41
R653 VDD.n193 VDD.n187 8629.41
R654 VDD.n206 VDD.n205 8629.41
R655 VDD.n208 VDD.n203 8629.41
R656 VDD.n226 VDD.n220 8629.41
R657 VDD.n229 VDD.n219 8629.41
R658 VDD.n242 VDD.n241 8629.41
R659 VDD.n244 VDD.n238 8629.41
R660 VDD.n259 VDD.n252 8629.41
R661 VDD.n256 VDD.n253 8629.41
R662 VDD.n53 VDD.n52 8629.41
R663 VDD.n55 VDD.n50 8629.41
R664 VDD.n36 VDD.n35 8629.41
R665 VDD.n38 VDD.n33 8629.41
R666 VDD.n19 VDD.n17 8629.41
R667 VDD.n22 VDD.n16 8629.41
R668 VDD.n8 VDD.n2 8629.41
R669 VDD.n8 VDD.n3 8629.41
R670 VDD.n6 VDD.n2 8629.41
R671 VDD.n6 VDD.n3 8629.41
R672 VDD.n276 VDD.n270 8629.41
R673 VDD.n276 VDD.n271 8629.41
R674 VDD.n274 VDD.n270 8629.41
R675 VDD.n274 VDD.n271 8629.41
R676 VDD.n8 VDD.t75 2459.29
R677 VDD.t76 VDD.n6 2459.29
R678 VDD.n276 VDD.t5 2459.29
R679 VDD.t2 VDD.n274 2459.29
R680 VDD.t75 VDD.n7 2298.92
R681 VDD.n7 VDD.t76 2298.92
R682 VDD.t5 VDD.n275 2298.92
R683 VDD.n275 VDD.t2 2298.92
R684 VDD.n189 VDD.n186 920.471
R685 VDD.n209 VDD.n202 920.471
R686 VDD.n225 VDD.n221 920.471
R687 VDD.n245 VDD.n237 920.471
R688 VDD.n255 VDD.n254 920.471
R689 VDD.n56 VDD.n49 920.471
R690 VDD.n39 VDD.n32 920.471
R691 VDD.n18 VDD.n15 920.471
R692 VDD.n5 VDD.n4 920.471
R693 VDD.n273 VDD.n272 920.471
R694 VDD.n195 VDD.n186 914.447
R695 VDD.n210 VDD.n209 914.447
R696 VDD.n221 VDD.n217 914.447
R697 VDD.n246 VDD.n245 914.447
R698 VDD.n254 VDD.n251 914.447
R699 VDD.n58 VDD.n56 914.447
R700 VDD.n41 VDD.n39 914.447
R701 VDD.n24 VDD.n15 914.447
R702 VDD.n4 VDD.n0 914.447
R703 VDD.n272 VDD.n268 914.447
R704 VDD.t68 VDD.n124 804.731
R705 VDD.n126 VDD.t68 751.692
R706 VDD.n98 VDD.t56 671.408
R707 VDD.n87 VDD.t47 671.408
R708 VDD VDD.t67 630.375
R709 VDD.n157 VDD.n156 602.456
R710 VDD.n179 VDD.n67 602.456
R711 VDD.n71 VDD.n70 585
R712 VDD.n73 VDD.n72 585
R713 VDD.n5 VDD.n1 480.764
R714 VDD.n273 VDD.n269 480.764
R715 VDD.n189 VDD.n184 480.764
R716 VDD.n202 VDD.n200 480.764
R717 VDD.n225 VDD.n224 480.764
R718 VDD.n239 VDD.n237 480.764
R719 VDD.n255 VDD.n250 480.764
R720 VDD.n49 VDD.n47 480.764
R721 VDD.n32 VDD.n30 480.764
R722 VDD.n18 VDD.n14 480.764
R723 VDD VDD.t70 458.724
R724 VDD.t67 VDD 458.724
R725 VDD.n119 VDD.t0 420.25
R726 VDD.n115 VDD.t71 388.656
R727 VDD.n150 VDD.t72 388.656
R728 VDD.n128 VDD.t69 388.656
R729 VDD.n101 VDD.t65 388.656
R730 VDD.n110 VDD.t66 388.656
R731 VDD.n75 VDD.t62 388.656
R732 VDD.n80 VDD.t63 388.656
R733 VDD.n197 VDD.n184 379.2
R734 VDD.n212 VDD.n200 379.2
R735 VDD.n224 VDD.n223 379.2
R736 VDD.n239 VDD.n236 379.2
R737 VDD.n263 VDD.n250 379.2
R738 VDD.n60 VDD.n47 379.2
R739 VDD.n43 VDD.n30 379.2
R740 VDD.n26 VDD.n14 379.2
R741 VDD.n10 VDD.n1 379.2
R742 VDD.n278 VDD.n269 379.2
R743 VDD VDD.t57 369.938
R744 VDD VDD.t77 369.938
R745 VDD.n104 VDD.n97 322.329
R746 VDD.n82 VDD.n78 322.329
R747 VDD.n161 VDD.n159 259.697
R748 VDD.n137 VDD.t78 255.905
R749 VDD.n142 VDD.t58 255.905
R750 VDD.n118 VDD.t1 255.905
R751 VDD.n158 VDD.t14 255.905
R752 VDD.n108 VDD.t34 254.475
R753 VDD.n133 VDD.t19 252.95
R754 VDD.n138 VDD.t54 252.95
R755 VDD.n143 VDD.t4 252.95
R756 VDD.n178 VDD.t30 252.95
R757 VDD.n157 VDD.t24 251.516
R758 VDD.n68 VDD.t74 250.724
R759 VDD.n66 VDD.t32 250.724
R760 VDD.t0 VDD.t3 248.599
R761 VDD.t57 VDD.t53 248.599
R762 VDD.t77 VDD.t18 248.599
R763 VDD.n173 VDD.t26 248.219
R764 VDD.n160 VDD.t12 248.219
R765 VDD.n119 VDD 221.964
R766 VDD.n126 VDD.t81 215.827
R767 VDD.n108 VDD.n107 213.119
R768 VDD.n148 VDD.n119 213.119
R769 VDD.n116 VDD.t80 210.964
R770 VDD.n102 VDD.t82 210.964
R771 VDD.n77 VDD.t79 210.964
R772 VDD.n168 VDD.n167 209.368
R773 VDD.t3 VDD 198.287
R774 VDD.t53 VDD 198.287
R775 VDD.t18 VDD 198.287
R776 VDD.n170 VDD.n169 183.673
R777 VDD VDD.t35 182.952
R778 VDD VDD.n168 182.952
R779 VDD.t37 VDD 182.952
R780 VDD.n72 VDD.n71 159.476
R781 VDD.n159 VDD.t50 157.014
R782 VDD.t73 VDD.t8 154.417
R783 VDD.t15 VDD.t13 147.703
R784 VDD.t48 VDD.t55 140.989
R785 VDD.t13 VDD.t11 140.989
R786 VDD.t29 VDD.t31 140.989
R787 VDD.t25 VDD.t73 140.989
R788 VDD.t46 VDD.t43 140.989
R789 VDD.n159 VDD.t40 137.079
R790 VDD.n107 VDD 125.883
R791 VDD.n169 VDD 125.883
R792 VDD.n97 VDD.t49 116.341
R793 VDD.n78 VDD.t44 116.341
R794 VDD.t55 VDD 112.457
R795 VDD.t11 VDD 112.457
R796 VDD VDD.t46 112.457
R797 VDD VDD.t59 109.1
R798 VDD.n11 VDD.n0 105.788
R799 VDD.n279 VDD.n268 105.788
R800 VDD.t64 VDD.t48 104.064
R801 VDD.t43 VDD.t61 104.064
R802 VDD.t27 VDD 102.385
R803 VDD.t33 VDD 99.0288
R804 VDD.n156 VDD.t16 96.1553
R805 VDD.n67 VDD.t21 96.1553
R806 VDD VDD.t20 92.315
R807 VDD.n71 VDD.t9 86.7743
R808 VDD.n107 VDD.t33 83.9228
R809 VDD.n168 VDD.t39 80.5659
R810 VDD.t35 VDD.t64 77.209
R811 VDD.t61 VDD.t37 77.209
R812 VDD.n72 VDD.t60 66.8398
R813 VDD.n196 VDD.n195 66.6358
R814 VDD.n211 VDD.n210 66.6358
R815 VDD.n218 VDD.n217 66.6358
R816 VDD.n247 VDD.n246 66.6358
R817 VDD.n262 VDD.n251 66.6358
R818 VDD.n59 VDD.n58 66.6358
R819 VDD.n42 VDD.n41 66.6358
R820 VDD.n25 VDD.n24 66.6358
R821 VDD.n10 VDD.n9 63.3551
R822 VDD.n278 VDD.n277 63.3551
R823 VDD.n156 VDD.t28 63.3219
R824 VDD.n67 VDD.t52 63.3219
R825 VDD VDD.t15 62.103
R826 VDD.n190 VDD.n189 61.6672
R827 VDD.n194 VDD.n193 61.6672
R828 VDD.n206 VDD.n202 61.6672
R829 VDD.n203 VDD.n201 61.6672
R830 VDD.n226 VDD.n225 61.6672
R831 VDD.n230 VDD.n229 61.6672
R832 VDD.n242 VDD.n237 61.6672
R833 VDD.n238 VDD.n234 61.6672
R834 VDD.n260 VDD.n259 61.6672
R835 VDD.n256 VDD.n255 61.6672
R836 VDD.n53 VDD.n49 61.6672
R837 VDD.n50 VDD.n48 61.6672
R838 VDD.n36 VDD.n32 61.6672
R839 VDD.n33 VDD.n31 61.6672
R840 VDD.n19 VDD.n18 61.6672
R841 VDD.n23 VDD.n22 61.6672
R842 VDD.n6 VDD.n5 61.6672
R843 VDD.n9 VDD.n8 61.6672
R844 VDD.n274 VDD.n273 61.6672
R845 VDD.n277 VDD.n276 61.6672
R846 VDD.n191 VDD.n190 60.9564
R847 VDD.n193 VDD.n192 60.9564
R848 VDD.n207 VDD.n206 60.9564
R849 VDD.n204 VDD.n203 60.9564
R850 VDD.n227 VDD.n226 60.9564
R851 VDD.n229 VDD.n228 60.9564
R852 VDD.n243 VDD.n242 60.9564
R853 VDD.n240 VDD.n238 60.9564
R854 VDD.n259 VDD.n258 60.9564
R855 VDD.n257 VDD.n256 60.9564
R856 VDD.n54 VDD.n53 60.9564
R857 VDD.n51 VDD.n50 60.9564
R858 VDD.n37 VDD.n36 60.9564
R859 VDD.n34 VDD.n33 60.9564
R860 VDD.n20 VDD.n19 60.9564
R861 VDD.n22 VDD.n21 60.9564
R862 VDD.n211 VDD.n201 60.6123
R863 VDD.n230 VDD.n218 60.6123
R864 VDD.n59 VDD.n48 60.6123
R865 VDD.n42 VDD.n31 60.6123
R866 VDD.n196 VDD.n185 59.4829
R867 VDD.n262 VDD.n261 59.4829
R868 VDD.n248 VDD.n247 58.7299
R869 VDD.n25 VDD.n13 58.7299
R870 VDD.t8 VDD 55.3892
R871 VDD.t51 VDD 52.0323
R872 VDD VDD.t39 45.3185
R873 VDD VDD.t23 41.9616
R874 VDD.n191 VDD.n187 38.5759
R875 VDD.n192 VDD.n188 38.5759
R876 VDD.n208 VDD.n207 38.5759
R877 VDD.n205 VDD.n204 38.5759
R878 VDD.n227 VDD.n219 38.5759
R879 VDD.n228 VDD.n220 38.5759
R880 VDD.n244 VDD.n243 38.5759
R881 VDD.n241 VDD.n240 38.5759
R882 VDD.n257 VDD.n252 38.5759
R883 VDD.n258 VDD.n253 38.5759
R884 VDD.n55 VDD.n54 38.5759
R885 VDD.n52 VDD.n51 38.5759
R886 VDD.n38 VDD.n37 38.5759
R887 VDD.n35 VDD.n34 38.5759
R888 VDD.n20 VDD.n16 38.5759
R889 VDD.n21 VDD.n17 38.5759
R890 VDD.n167 VDD.n89 34.6358
R891 VDD.n167 VDD.n90 34.6358
R892 VDD.n172 VDD.n171 34.6358
R893 VDD.n169 VDD 28.5341
R894 VDD.n97 VDD.t36 28.4453
R895 VDD.n78 VDD.t38 28.4453
R896 VDD.n174 VDD.n173 28.3534
R897 VDD.n171 VDD.n170 25.6953
R898 VDD.n137 VDD.n122 25.224
R899 VDD.n133 VDD.n122 25.224
R900 VDD.n142 VDD.n121 25.224
R901 VDD.n138 VDD.n121 25.224
R902 VDD.n144 VDD.n118 25.224
R903 VDD.n144 VDD.n143 25.224
R904 VDD.n162 VDD.n158 25.224
R905 VDD.n108 VDD.n92 23.7181
R906 VDD VDD.n98 23.252
R907 VDD.n157 VDD.n92 21.4593
R908 VDD.n138 VDD.n137 20.3299
R909 VDD.n143 VDD.n142 20.3299
R910 VDD.t20 VDD.t29 20.1418
R911 VDD.n179 VDD.n66 19.9534
R912 VDD.n178 VDD.n177 19.8181
R913 VDD.n148 VDD.n118 17.3181
R914 VDD.n161 VDD.n160 17.3181
R915 VDD.n158 VDD.n157 16.5652
R916 VDD.n162 VDD.n161 16.5652
R917 VDD.n133 VDD.n132 15.8123
R918 VDD.n149 VDD.n148 14.2735
R919 VDD.n109 VDD.n108 14.2735
R920 VDD.n171 VDD.n87 13.9299
R921 VDD.n179 VDD.n178 13.5534
R922 VDD.n114 VDD.n113 11.4366
R923 VDD.n198 VDD.n197 11.3235
R924 VDD.n213 VDD.n212 11.3235
R925 VDD.n223 VDD.n222 11.3235
R926 VDD.n236 VDD.n235 11.3235
R927 VDD.n264 VDD.n263 11.3235
R928 VDD.n61 VDD.n60 11.3235
R929 VDD.n44 VDD.n43 11.3235
R930 VDD.n27 VDD.n26 11.3235
R931 VDD.n170 VDD.n88 11.2937
R932 VDD.n154 VDD.n153 11.2737
R933 VDD.t23 VDD.t27 10.0712
R934 VDD.n128 VDD.n125 9.60526
R935 VDD.n115 VDD.n114 9.60526
R936 VDD.n80 VDD.n79 9.60526
R937 VDD.n117 VDD.n93 9.3005
R938 VDD.n152 VDD.n151 9.3005
R939 VDD.n149 VDD.n94 9.3005
R940 VDD.n148 VDD.n147 9.3005
R941 VDD.n143 VDD.n120 9.3005
R942 VDD.n139 VDD.n138 9.3005
R943 VDD.n134 VDD.n133 9.3005
R944 VDD.n130 VDD.n129 9.3005
R945 VDD.n135 VDD.n122 9.3005
R946 VDD.n137 VDD.n136 9.3005
R947 VDD.n140 VDD.n121 9.3005
R948 VDD.n142 VDD.n141 9.3005
R949 VDD.n145 VDD.n144 9.3005
R950 VDD.n146 VDD.n118 9.3005
R951 VDD.n175 VDD.n174 9.3005
R952 VDD.n180 VDD.n179 9.3005
R953 VDD.n164 VDD.n89 9.3005
R954 VDD.n157 VDD.n155 9.3005
R955 VDD.n108 VDD.n106 9.3005
R956 VDD.n100 VDD.n99 9.3005
R957 VDD.n103 VDD.n95 9.3005
R958 VDD.n112 VDD.n111 9.3005
R959 VDD.n109 VDD.n96 9.3005
R960 VDD.n105 VDD.n92 9.3005
R961 VDD.n158 VDD.n91 9.3005
R962 VDD.n163 VDD.n162 9.3005
R963 VDD.n167 VDD.n166 9.3005
R964 VDD.n165 VDD.n90 9.3005
R965 VDD.n178 VDD.n65 9.3005
R966 VDD.n177 VDD.n176 9.3005
R967 VDD.n172 VDD.n69 9.3005
R968 VDD.n171 VDD.n74 9.3005
R969 VDD.n86 VDD.n85 9.3005
R970 VDD.n84 VDD.n83 9.3005
R971 VDD.n81 VDD.n76 9.3005
R972 VDD.n28 VDD.n13 8.23557
R973 VDD.n12 VDD.n11 7.54844
R974 VDD.n280 VDD.n279 7.54407
R975 VDD.n185 VDD.n183 6.88686
R976 VDD.n73 VDD.n70 6.8005
R977 VDD.n132 VDD.n124 6.48583
R978 VDD.n195 VDD.n194 6.02403
R979 VDD.n246 VDD.n234 6.02403
R980 VDD.n260 VDD.n251 6.02403
R981 VDD.n24 VDD.n23 6.02403
R982 VDD.n9 VDD.n0 6.02403
R983 VDD.n277 VDD.n268 6.02403
R984 VDD.n127 VDD.n126 5.8885
R985 VDD.n11 VDD.n10 5.18145
R986 VDD.n279 VDD.n278 5.18145
R987 VDD.n201 VDD.n64 4.89462
R988 VDD.n231 VDD.n217 4.89462
R989 VDD.n57 VDD.n48 4.89462
R990 VDD.n41 VDD.n40 4.89462
R991 VDD.n151 VDD.n117 4.67352
R992 VDD.n132 VDD.n131 4.62124
R993 VDD.n129 VDD.n128 4.36875
R994 VDD.n151 VDD.n150 4.36875
R995 VDD.n111 VDD.n110 4.36875
R996 VDD.n81 VDD.n80 4.36875
R997 VDD.t31 VDD.t51 3.35739
R998 VDD.t59 VDD.t25 3.35739
R999 VDD.n183 VDD 3.29986
R1000 VDD.n215 VDD.n64 3.25464
R1001 VDD.n249 VDD.n248 3.24308
R1002 VDD.n57 VDD.n46 3.23917
R1003 VDD.n232 VDD.n231 3.23136
R1004 VDD.n40 VDD.n29 3.23136
R1005 VDD.n261 VDD.n63 3.22655
R1006 VDD.n129 VDD.n127 3.2005
R1007 VDD.n187 VDD.n186 2.84665
R1008 VDD.n188 VDD.n184 2.84665
R1009 VDD.n209 VDD.n208 2.84665
R1010 VDD.n205 VDD.n200 2.84665
R1011 VDD.n221 VDD.n219 2.84665
R1012 VDD.n224 VDD.n220 2.84665
R1013 VDD.n245 VDD.n244 2.84665
R1014 VDD.n241 VDD.n239 2.84665
R1015 VDD.n254 VDD.n252 2.84665
R1016 VDD.n253 VDD.n250 2.84665
R1017 VDD.n56 VDD.n55 2.84665
R1018 VDD.n52 VDD.n47 2.84665
R1019 VDD.n39 VDD.n38 2.84665
R1020 VDD.n35 VDD.n30 2.84665
R1021 VDD.n16 VDD.n15 2.84665
R1022 VDD.n17 VDD.n14 2.84665
R1023 VDD.n3 VDD.n1 2.84665
R1024 VDD.n7 VDD.n3 2.84665
R1025 VDD.n4 VDD.n2 2.84665
R1026 VDD.n7 VDD.n2 2.84665
R1027 VDD.n271 VDD.n269 2.84665
R1028 VDD.n275 VDD.n271 2.84665
R1029 VDD.n272 VDD.n270 2.84665
R1030 VDD.n275 VDD.n270 2.84665
R1031 VDD.n127 VDD.n124 2.8165
R1032 VDD.n104 VDD.n103 2.54018
R1033 VDD.n83 VDD.n82 2.54018
R1034 VDD.n117 VDD.n116 2.33701
R1035 VDD.n103 VDD.n102 2.33701
R1036 VDD.n83 VDD.n77 2.33701
R1037 VDD.n197 VDD.n196 2.28169
R1038 VDD.n212 VDD.n211 2.28169
R1039 VDD.n223 VDD.n218 2.28169
R1040 VDD.n247 VDD.n236 2.28169
R1041 VDD.n263 VDD.n262 2.28169
R1042 VDD.n60 VDD.n59 2.28169
R1043 VDD.n43 VDD.n42 2.28169
R1044 VDD.n26 VDD.n25 2.28169
R1045 VDD.n233 VDD.n232 2.13544
R1046 VDD.n111 VDD.n104 2.13383
R1047 VDD.n82 VDD.n81 2.13383
R1048 VDD.n267 VDD.n12 2.06883
R1049 VDD.n116 VDD.n115 2.03225
R1050 VDD.n102 VDD.n101 2.03225
R1051 VDD.n77 VDD.n75 2.03225
R1052 VDD.n249 VDD.n233 1.95379
R1053 VDD.n248 VDD.n234 1.88285
R1054 VDD.n23 VDD.n13 1.88285
R1055 VDD.n182 VDD.n181 1.753
R1056 VDD VDD.n182 1.64258
R1057 VDD.n90 VDD.n66 1.50638
R1058 VDD.n174 VDD.n73 1.4005
R1059 VDD.n100 VDD.n98 1.37193
R1060 VDD.n87 VDD.n86 1.37193
R1061 VDD.n280 VDD.n267 1.33758
R1062 VDD.n214 VDD.n213 1.143
R1063 VDD.n222 VDD.n216 1.143
R1064 VDD.n62 VDD.n61 1.143
R1065 VDD.n45 VDD.n44 1.143
R1066 VDD.n199 VDD.n198 1.13925
R1067 VDD.n265 VDD.n264 1.13925
R1068 VDD.n235 VDD.n233 1.13675
R1069 VDD.n28 VDD.n27 1.13675
R1070 VDD.n194 VDD.n185 1.12991
R1071 VDD.n210 VDD.n64 1.12991
R1072 VDD.n231 VDD.n230 1.12991
R1073 VDD.n261 VDD.n260 1.12991
R1074 VDD.n58 VDD.n57 1.12991
R1075 VDD.n40 VDD.n31 1.12991
R1076 VDD.n123 VDD 1.06099
R1077 VDD.n46 VDD.n45 0.862816
R1078 VDD.n214 VDD.n199 0.854667
R1079 VDD.n29 VDD.n28 0.770881
R1080 VDD.n160 VDD.n89 0.753441
R1081 VDD.n173 VDD.n172 0.753441
R1082 VDD.n63 VDD.n62 0.747859
R1083 VDD.n267 VDD.n266 0.704667
R1084 VDD.n70 VDD.n68 0.6005
R1085 VDD.n216 VDD.n215 0.588641
R1086 VDD.n265 VDD.n249 0.518882
R1087 VDD.n182 VDD 0.460219
R1088 VDD.n177 VDD.n68 0.4005
R1089 VDD.n45 VDD.n29 0.392323
R1090 VDD.n62 VDD.n46 0.360318
R1091 VDD.n150 VDD.n149 0.305262
R1092 VDD.n101 VDD.n100 0.305262
R1093 VDD.n110 VDD.n109 0.305262
R1094 VDD.n86 VDD.n75 0.305262
R1095 VDD.t45 VDD.n191 0.27666
R1096 VDD.n192 VDD.t45 0.27666
R1097 VDD.n207 VDD.t17 0.27666
R1098 VDD.n204 VDD.t17 0.27666
R1099 VDD.t42 VDD.n227 0.27666
R1100 VDD.n228 VDD.t42 0.27666
R1101 VDD.n243 VDD.t10 0.27666
R1102 VDD.n240 VDD.t10 0.27666
R1103 VDD.t6 VDD.n257 0.27666
R1104 VDD.n258 VDD.t6 0.27666
R1105 VDD.n54 VDD.t7 0.27666
R1106 VDD.n51 VDD.t7 0.27666
R1107 VDD.n37 VDD.t41 0.27666
R1108 VDD.n34 VDD.t41 0.27666
R1109 VDD.t22 VDD.n20 0.27666
R1110 VDD.n21 VDD.t22 0.27666
R1111 VDD.n215 VDD.n214 0.268128
R1112 VDD.n232 VDD.n216 0.223986
R1113 VDD.n199 VDD.n183 0.202423
R1114 VDD.n131 VDD.n130 0.180304
R1115 VDD.n131 VDD 0.120408
R1116 VDD.n114 VDD.n93 0.120292
R1117 VDD.n152 VDD.n94 0.120292
R1118 VDD.n146 VDD.n145 0.120292
R1119 VDD.n145 VDD.n120 0.120292
R1120 VDD.n141 VDD.n140 0.120292
R1121 VDD.n140 VDD.n139 0.120292
R1122 VDD.n136 VDD.n135 0.120292
R1123 VDD.n135 VDD.n134 0.120292
R1124 VDD.n130 VDD.n125 0.120292
R1125 VDD.n99 VDD.n95 0.120292
R1126 VDD.n112 VDD.n96 0.120292
R1127 VDD.n163 VDD.n91 0.120292
R1128 VDD.n164 VDD.n163 0.120292
R1129 VDD.n180 VDD.n65 0.120292
R1130 VDD.n176 VDD.n175 0.120292
R1131 VDD.n175 VDD.n69 0.120292
R1132 VDD.n85 VDD.n84 0.120292
R1133 VDD.n84 VDD.n76 0.120292
R1134 VDD.n79 VDD.n76 0.120292
R1135 VDD.n153 VDD.n93 0.11899
R1136 VDD.n266 VDD.n63 0.1125
R1137 VDD.n99 VDD 0.0981562
R1138 VDD.n154 VDD 0.0955521
R1139 VDD.n113 VDD.n95 0.0916458
R1140 VDD.n198 VDD 0.06425
R1141 VDD.n213 VDD 0.06425
R1142 VDD.n222 VDD 0.06425
R1143 VDD.n235 VDD 0.06425
R1144 VDD.n264 VDD 0.06425
R1145 VDD.n61 VDD 0.06425
R1146 VDD.n44 VDD 0.06425
R1147 VDD.n27 VDD 0.06425
R1148 VDD VDD.n280 0.06425
R1149 VDD.n147 VDD 0.0603958
R1150 VDD VDD.n146 0.0603958
R1151 VDD.n141 VDD 0.0603958
R1152 VDD.n136 VDD 0.0603958
R1153 VDD.n106 VDD 0.0603958
R1154 VDD VDD.n105 0.0603958
R1155 VDD VDD.n91 0.0603958
R1156 VDD.n166 VDD 0.0603958
R1157 VDD VDD.n165 0.0603958
R1158 VDD.n176 VDD 0.0603958
R1159 VDD.n85 VDD 0.0603958
R1160 VDD.n12 VDD 0.059875
R1161 VDD.n88 VDD 0.0590938
R1162 VDD.n266 VDD.n265 0.054
R1163 VDD.n181 VDD 0.0525833
R1164 VDD.n181 VDD.n180 0.0460729
R1165 VDD.n106 VDD 0.0382604
R1166 VDD VDD.n123 0.0369583
R1167 VDD.n147 VDD 0.03175
R1168 VDD.n166 VDD 0.03175
R1169 VDD.n113 VDD.n112 0.0291458
R1170 VDD VDD.n94 0.0226354
R1171 VDD VDD.n120 0.0226354
R1172 VDD.n139 VDD 0.0226354
R1173 VDD.n134 VDD 0.0226354
R1174 VDD.n125 VDD 0.0226354
R1175 VDD VDD.n96 0.0226354
R1176 VDD.n105 VDD 0.0226354
R1177 VDD.n155 VDD 0.0226354
R1178 VDD VDD.n164 0.0226354
R1179 VDD.n165 VDD 0.0226354
R1180 VDD VDD.n65 0.0226354
R1181 VDD VDD.n69 0.0226354
R1182 VDD VDD.n74 0.0226354
R1183 VDD.n79 VDD 0.0226354
R1184 VDD.n155 VDD.n154 0.00310417
R1185 VDD.n153 VDD.n152 0.00180208
R1186 VDD.n123 VDD 0.00180208
R1187 VDD.n88 VDD.n74 0.00180208
R1188 x3.GN1.n2 x3.GN1.t9 377.486
R1189 x3.GN1.n3 x3.GN1.t2 377.486
R1190 x3.GN1.n2 x3.GN1.t7 374.202
R1191 x3.GN1.n3 x3.GN1.t3 374.202
R1192 x3.GN1.n10 x3.GN1.t0 339.418
R1193 x3.GN1.n1 x3.GN1.t1 274.06
R1194 x3.GN1.n7 x3.GN1.t8 212.081
R1195 x3.GN1.n6 x3.GN1.t6 212.081
R1196 x3.GN1.n8 x3.GN1.n7 182.673
R1197 x3.GN1.n7 x3.GN1.t5 139.78
R1198 x3.GN1.n6 x3.GN1.t4 139.78
R1199 x3.GN1.n7 x3.GN1.n6 61.346
R1200 x3.GN1.n5 x3.GN1.n8 15.8606
R1201 x3.GN1 x3.GN1.n9 13.8044
R1202 x3.GN1.n0 x3.GN1.n4 13.4101
R1203 x3.GN1.n0 x3.GN1 11.6184
R1204 x3.GN1.n4 x3.GN1 11.6184
R1205 x3.GN1 x3.GN1.n1 11.0989
R1206 x3.GN1.n9 x3.GN1.n5 6.94768
R1207 x3.GN1 x3.GN1.n0 6.73859
R1208 x3.GN1.n11 x3.GN1 6.6565
R1209 x3.GN1.n8 x3.GN1 6.4005
R1210 x3.GN1.n1 x3.GN1 6.1445
R1211 x3.GN1.n0 x3.GN1 5.13959
R1212 x3.GN1.n4 x3.GN1 4.55738
R1213 x3.GN1.n11 x3.GN1.n10 4.0914
R1214 x3.GN1 x3.GN1.n11 3.61789
R1215 x3.GN1.n9 x3.GN1 3.26325
R1216 x3.GN1.n1 x3.GN1 2.86947
R1217 x3.GN1 x3.GN1.n3 2.04102
R1218 x3.GN1 x3.GN1.n2 2.04102
R1219 x3.GN1.n10 x3.GN1 1.74382
R1220 x3.GN1.n5 x3.GN1 1.47326
R1221 A5.n1 A5.t0 26.3998
R1222 A5.n1 A5.t3 23.5483
R1223 A5.n0 A5.t2 12.7127
R1224 A5.n0 A5.t1 10.8578
R1225 A5.n2 A5.n1 3.12177
R1226 A5.n2 A5.n0 1.81453
R1227 A5.n3 A5.n2 1.1255
R1228 A5.n3 A5 0.21549
R1229 A5 A5.n3 0.0655
R1230 x3.GN4.n3 x3.GN4.t3 377.486
R1231 x3.GN4.n1 x3.GN4.t6 377.486
R1232 x3.GN4.n3 x3.GN4.t5 374.202
R1233 x3.GN4.n1 x3.GN4.t9 374.202
R1234 x3.GN4.n9 x3.GN4.t0 339.418
R1235 x3.GN4.n0 x3.GN4.t1 274.06
R1236 x3.GN4.n6 x3.GN4.t4 212.081
R1237 x3.GN4.n5 x3.GN4.t8 212.081
R1238 x3.GN4.n7 x3.GN4.n6 184.977
R1239 x3.GN4.n6 x3.GN4.t2 139.78
R1240 x3.GN4.n5 x3.GN4.t7 139.78
R1241 x3.GN4.n6 x3.GN4.n5 61.346
R1242 x3.GN4.n8 x3.GN4 18.2601
R1243 x3.GN4 x3.GN4.n7 13.8193
R1244 x3.GN4 x3.GN4.n4 11.7568
R1245 x3.GN4.n4 x3.GN4.n2 11.6628
R1246 x3.GN4 x3.GN4.n0 11.2645
R1247 x3.GN4 x3.GN4.n8 8.9605
R1248 x3.GN4.n8 x3.GN4 8.4485
R1249 x3.GN4.n2 x3.GN4 8.19806
R1250 x3.GN4.n10 x3.GN4 6.6565
R1251 x3.GN4.n0 x3.GN4 6.1445
R1252 x3.GN4.n4 x3.GN4 5.8185
R1253 x3.GN4.n2 x3.GN4 4.58237
R1254 x3.GN4.n7 x3.GN4 4.0965
R1255 x3.GN4.n10 x3.GN4.n9 4.0914
R1256 x3.GN4 x3.GN4.n10 3.61789
R1257 x3.GN4.n0 x3.GN4 2.86947
R1258 x3.GN4 x3.GN4.n1 2.04102
R1259 x3.GN4 x3.GN4.n3 2.04102
R1260 x3.GN4.n9 x3.GN4 1.74382
R1261 x3.GP4.n3 x3.GP4.t7 450.938
R1262 x3.GP4.n2 x3.GP4.t4 450.938
R1263 x3.GP4.n3 x3.GP4.t5 445.666
R1264 x3.GP4.n2 x3.GP4.t6 445.666
R1265 x1.x14.Y x3.GP4.n7 203.923
R1266 x3.GP4.n1 x3.GP4.n0 101.49
R1267 x3.GP4.n7 x3.GP4.t0 26.5955
R1268 x3.GP4.n7 x3.GP4.t1 26.5955
R1269 x3.GP4.n0 x3.GP4.t2 24.9236
R1270 x3.GP4.n0 x3.GP4.t3 24.9236
R1271 x3.GP4.n4 x3.x4.GP 11.0619
R1272 x3.GP4.n6 x1.x14.Y 10.7525
R1273 x1.gpo3 x3.GP4.n4 9.34192
R1274 x3.GP4.n5 x1.gpo3 7.73829
R1275 x3.GP4.n6 x1.x14.Y 6.6565
R1276 x3.GP4.n4 x2.x4.GP 5.84951
R1277 x1.x14.Y x3.GP4.n6 5.04292
R1278 x2.x4.GP x3.GP4.n3 2.95993
R1279 x3.x4.GP x3.GP4.n2 2.95993
R1280 x3.GP4.n1 x1.x14.Y 1.93989
R1281 x1.x14.Y x3.GP4.n5 1.5365
R1282 x3.GP4.n5 x3.GP4.n1 1.0245
R1283 select0.n5 select0.t3 327.99
R1284 select0.n9 select0.t2 293.969
R1285 select0.n3 select0.t6 261.887
R1286 select0.n1 select0.t1 212.081
R1287 select0.n0 select0.t0 212.081
R1288 select0.n5 select0.t5 199.457
R1289 select0.n2 select0.n1 183.185
R1290 select0.n3 select0.t4 155.847
R1291 select0 select0.n9 154.065
R1292 select0.n6 select0.n5 152
R1293 select0.n4 select0.n3 152
R1294 select0.n1 select0.t9 139.78
R1295 select0.n0 select0.t8 139.78
R1296 select0.n9 select0.t7 138.338
R1297 select0.n1 select0.n0 61.346
R1298 select0.n10 select0 13.4199
R1299 select0.n8 select0.n4 11.9062
R1300 select0.n11 select0.n8 11.7395
R1301 select0.n12 select0.n11 11.5949
R1302 select0.n12 select0.n2 9.68118
R1303 select0.n7 select0 9.17383
R1304 select0.n2 select0 5.8885
R1305 select0.n10 select0 5.57469
R1306 select0.n8 select0.n7 4.6505
R1307 select0.n11 select0.n10 4.6505
R1308 select0.n7 select0.n6 2.98717
R1309 select0.n6 select0 2.34717
R1310 select0.n4 select0 2.07109
R1311 select0 select0.n12 0.559212
R1312 x3.GP1.n4 x3.GP1.t5 450.938
R1313 x3.GP1.n3 x3.GP1.t7 450.938
R1314 x3.GP1.n4 x3.GP1.t4 445.666
R1315 x3.GP1.n3 x3.GP1.t6 445.666
R1316 x3.GP1.n7 x3.GP1.n6 195.832
R1317 x3.GP1.n1 x3.GP1.n0 101.49
R1318 x3.GP1.n6 x3.GP1.t1 26.5955
R1319 x3.GP1.n6 x3.GP1.t0 26.5955
R1320 x3.GP1.n0 x3.GP1.t3 24.9236
R1321 x3.GP1.n0 x3.GP1.t2 24.9236
R1322 x3.GP1.n5 x3.x1.GP 13.3282
R1323 x3.GP1.n7 x1.gpo0 11.8923
R1324 x3.GP1.n2 x1.x11.Y 10.7525
R1325 x1.x11.Y x3.GP1.n7 8.09215
R1326 x3.GP1.n2 x1.x11.Y 6.6565
R1327 x1.gpo0 x3.GP1.n5 5.46644
R1328 x3.GP1.n5 x2.GP1 5.31412
R1329 x1.x11.Y x3.GP1.n2 5.04292
R1330 x2.GP1 x3.GP1.n4 3.18415
R1331 x3.x1.GP x3.GP1.n3 2.90754
R1332 x1.x11.Y x3.GP1.n1 2.5605
R1333 x3.GP1.n1 x1.x11.Y 1.93989
R1334 A1.n1 A1.t0 26.3998
R1335 A1.n1 A1.t1 23.5483
R1336 A1.n0 A1.t2 12.7127
R1337 A1.n0 A1.t3 10.8578
R1338 A1.n2 A1.n1 3.12177
R1339 A1.n2 A1.n0 1.81453
R1340 A1.n3 A1.n2 1.1255
R1341 A1.n3 A1 0.21549
R1342 A1 A1.n3 0.0655
R1343 A2.n1 A2.t0 26.3998
R1344 A2.n1 A2.t3 23.5483
R1345 A2.n0 A2.t1 12.7127
R1346 A2.n0 A2.t2 10.8578
R1347 A2.n2 A2.n1 3.12177
R1348 A2.n2 A2.n0 1.81453
R1349 A2.n3 A2.n2 1.1255
R1350 A2.n3 A2 0.219402
R1351 A2 A2.n3 0.0655
R1352 A4.n1 A4.t2 26.3998
R1353 A4.n1 A4.t3 23.5483
R1354 A4.n0 A4.t1 12.7127
R1355 A4.n0 A4.t0 10.8578
R1356 A4.n2 A4.n1 3.12177
R1357 A4.n2 A4.n0 1.81453
R1358 A4.n3 A4.n2 1.1255
R1359 A4 A4.n3 0.203263
R1360 A4.n3 A4 0.0655
R1361 A7.n1 A7.t2 26.3998
R1362 A7.n1 A7.t3 23.5483
R1363 A7.n0 A7.t1 12.7127
R1364 A7.n0 A7.t0 10.8578
R1365 A7.n2 A7.n1 3.12177
R1366 A7.n2 A7.n0 1.81453
R1367 A7.n3 A7.n2 1.1255
R1368 A7.n3 A7 0.210543
R1369 A7 A7.n3 0.0655
R1370 A3.n1 A3.t3 26.3998
R1371 A3.n1 A3.t2 23.5483
R1372 A3.n0 A3.t1 12.7127
R1373 A3.n0 A3.t0 10.8578
R1374 A3.n2 A3.n1 3.12177
R1375 A3.n2 A3.n0 1.81453
R1376 A3.n3 A3.n2 1.1255
R1377 A3.n3 A3 0.210543
R1378 A3 A3.n3 0.0655
R1379 A6.n1 A6.t3 26.3998
R1380 A6.n1 A6.t0 23.5483
R1381 A6.n0 A6.t2 12.7127
R1382 A6.n0 A6.t1 10.8578
R1383 A6.n2 A6.n1 3.12177
R1384 A6.n2 A6.n0 1.81453
R1385 A6.n3 A6.n2 1.1255
R1386 A6.n3 A6 0.219402
R1387 A6 A6.n3 0.0655
R1388 A8.n1 A8.t3 26.3998
R1389 A8.n1 A8.t2 23.5483
R1390 A8.n0 A8.t1 12.7127
R1391 A8.n0 A8.t0 10.8578
R1392 A8.n2 A8.n1 3.12177
R1393 A8.n2 A8.n0 1.81453
R1394 A8.n3 A8.n2 1.1255
R1395 A8 A8.n3 0.203263
R1396 A8.n3 A8 0.0655
R1397 x3.GP2.n4 x3.GP2.t6 450.938
R1398 x3.GP2.n3 x3.GP2.t7 450.938
R1399 x3.GP2.n4 x3.GP2.t4 445.666
R1400 x3.GP2.n3 x3.GP2.t5 445.666
R1401 x3.GP2.n7 x3.GP2.n6 195.958
R1402 x3.GP2.n1 x3.GP2.n0 101.49
R1403 x3.GP2.n6 x3.GP2.t1 26.5955
R1404 x3.GP2.n6 x3.GP2.t0 26.5955
R1405 x3.GP2.n0 x3.GP2.t3 24.9236
R1406 x3.GP2.n0 x3.GP2.t2 24.9236
R1407 x3.GP2.n5 x3.x2.GP 14.964
R1408 x3.GP2.n7 x1.gpo1 11.8408
R1409 x3.GP2.n2 x1.x12.Y 10.7525
R1410 x1.gpo1 x3.GP2.n5 8.86265
R1411 x1.x12.Y x3.GP2.n7 7.96524
R1412 x3.GP2.n2 x1.x12.Y 6.6565
R1413 x3.GP2.n5 x2.x2.GP 5.75481
R1414 x1.x12.Y x3.GP2.n2 5.04292
R1415 x2.x2.GP x3.GP2.n4 2.94361
R1416 x3.x2.GP x3.GP2.n3 2.94361
R1417 x1.x12.Y x3.GP2.n1 2.5605
R1418 x3.GP2.n1 x1.x12.Y 1.93989
C0 x3.GN1 A3 0.131584f
C1 VDD A4 1.56602f
C2 a_5645_6637# x3.GN4 0.003645f
C3 x4.A A8 4.51511f
C4 x3.GN3 a_5699_7287# 1.07e-20
C5 a_5645_6637# select1 0.127717f
C6 a_5699_7287# x3.GN4 0.001562f
C7 x3.GN1 x1.nSEL0 0.002613f
C8 a_5699_7287# select1 8.84e-19
C9 a_5645_6461# select0 0.086353f
C10 x3.GN1 a_5645_5909# 0.012357f
C11 VDD a_5645_7149# 0.217381f
C12 a_5645_6085# x5.GN 3.26e-19
C13 a_5645_6085# x3.GN3 0.048646f
C14 A3 VDD 1.61205f
C15 x5.GN a_5671_6037# 1.08e-19
C16 x3.GN3 a_5671_6037# 5.17e-20
C17 a_5645_6085# select1 0.254026f
C18 x3.GN1 a_5645_6461# 7.95e-20
C19 a_5645_6461# a_5671_6589# 0.004764f
C20 VDD x1.nSEL0 0.386805f
C21 x4.A select2 4.96806f
C22 x3.GN2 x4.A 0.429477f
C23 VDD a_5645_5909# 0.162117f
C24 x4.A x5.A 2.05508f
C25 x4.A x3.GP3 0.358391f
C26 a_5645_6637# select0 0.279858f
C27 A4 select2 6.76e-20
C28 m2_5776_5494# x5.GN 4e-19
C29 VDD a_5645_6461# 0.171399f
C30 x3.GN2 A4 6.05e-19
C31 x5.GN Z 0.820847f
C32 A4 x5.A 4.5151f
C33 a_5699_7287# select0 1.4e-19
C34 m2_5776_5494# select1 0.183786f
C35 A4 x3.GP3 0.162086f
C36 a_5645_5493# m2_5776_5494# 0.01297f
C37 x3.GN4 Z 9.07e-20
C38 x3.GN1 a_5645_6637# 1.69e-20
C39 x3.GN2 a_5645_7149# 7.58e-21
C40 a_5645_6085# select0 0.143958f
C41 x1.nSEL0 x1.nSEL1 0.352716f
C42 A3 select2 2.39e-19
C43 A3 x3.GN2 0.007138f
C44 x1.nSEL1 a_5645_5909# 0.073392f
C45 A3 x5.A 4.5214f
C46 A3 x3.GP3 3.96087f
C47 x1.nSEL0 select2 0.131256f
C48 x3.GN3 x5.GN 1.63e-19
C49 x1.nSEL0 x3.GN2 0.154394f
C50 select2 a_5645_5909# 8.66e-20
C51 a_5645_6637# VDD 0.262163f
C52 x3.GN1 a_5645_6085# 1.45e-19
C53 x3.GN2 a_5645_5909# 0.106139f
C54 x5.GN x3.GN4 9.02e-19
C55 x3.GN3 x3.GN4 0.195262f
C56 a_5645_6461# x1.nSEL1 7.84e-19
C57 select1 x5.GN 0.140519f
C58 x3.GN3 select1 0.272271f
C59 a_5645_5493# x5.GN 0.001336f
C60 x3.GN1 a_5671_6037# 1.22e-20
C61 VDD a_5699_7287# 8.97e-19
C62 select1 x3.GN4 0.059776f
C63 a_5645_5493# select1 0.02803f
C64 a_5645_6461# select2 0.009143f
C65 x3.GN2 a_5645_6461# 1.61e-19
C66 m2_5776_5494# select0 0.130999f
C67 x3.GN3 A7 3.80783f
C68 A4 x4.A 0.003925f
C69 VDD a_5645_6085# 0.193284f
C70 a_5645_6461# x3.GP3 0.001353f
C71 x3.GN4 A7 0.180503f
C72 VDD a_5671_6037# 4.32e-19
C73 x3.GN1 m2_5776_5494# 0.06935f
C74 x3.GN1 Z 4.27e-20
C75 A5 x3.GN3 2.86e-19
C76 a_5645_6637# x1.nSEL1 1.59e-19
C77 A3 x4.A 1.64e-20
C78 A5 x3.GN4 0.005885f
C79 x5.GN select0 0.131913f
C80 x3.GN3 select0 0.254198f
C81 a_5645_6637# x3.GN2 1.03e-19
C82 x3.GN4 select0 0.218342f
C83 m2_5776_5494# VDD 0.139797f
C84 select1 select0 1.85585f
C85 a_5645_5493# select0 0.048888f
C86 A3 A4 2.08862f
C87 x3.GN3 A2 0.137879f
C88 a_5645_6637# x3.GP3 4.69e-19
C89 x3.GN2 a_5699_7287# 8.14e-21
C90 VDD Z 5.306779f
C91 a_5645_6085# x1.nSEL1 0.041068f
C92 A6 x3.GN3 0.156179f
C93 x3.GN4 A2 1.76e-19
C94 A6 x3.GN4 1.76e-19
C95 x3.GN1 x5.GN 0.645008f
C96 x3.GN1 x3.GN3 0.089083f
C97 x1.nSEL1 a_5671_6037# 9.57e-19
C98 x5.GN a_5671_6589# 9.76e-20
C99 x3.GN3 a_5671_6589# 0.001073f
C100 x3.GN1 x3.GN4 0.14554f
C101 x3.GN4 a_5671_6589# 3.22e-19
C102 a_5645_6085# select2 1.67e-19
C103 a_5645_6085# x3.GN2 0.016995f
C104 x3.GN1 select1 0.312176f
C105 a_5645_5493# x3.GN1 0.128677f
C106 x3.GN2 a_5671_6037# 0.002395f
C107 A6 A7 1.81997f
C108 a_5699_5631# x5.GN 1.95e-19
C109 VDD x5.GN 3.62413f
C110 VDD x3.GN3 0.768845f
C111 VDD x3.GN4 1.35712f
C112 a_5645_5493# a_5699_5631# 0.006584f
C113 m2_5776_5494# x1.nSEL1 0.00815f
C114 VDD select1 2.65613f
C115 a_5645_5493# VDD 0.21052f
C116 A5 A6 1.81909f
C117 x3.GN3 A8 0.006957f
C118 x1.nSEL0 a_5645_5909# 0.03096f
C119 m2_5776_5494# select2 4.4e-19
C120 A5 x3.GN1 3.85245f
C121 select2 Z 0.76903f
C122 x3.GN4 A8 3.84613f
C123 x3.GN2 Z 9.36e-20
C124 VDD A7 1.61205f
C125 x5.A Z 4.51579f
C126 x3.GP3 Z 2.44e-19
C127 x3.GN1 select0 0.020289f
C128 x1.nSEL0 a_5645_6461# 1.91e-20
C129 a_5671_6589# select0 0.001558f
C130 x1.nSEL1 x5.GN 0.10521f
C131 x3.GN3 x1.nSEL1 0.012418f
C132 x3.GN1 A2 0.135398f
C133 A7 A8 2.08862f
C134 A5 VDD 1.60179f
C135 x3.GN1 A6 3.66e-20
C136 select1 x1.nSEL1 0.275603f
C137 a_5645_5493# x1.nSEL1 0.193944f
C138 select2 x5.GN 3.99214f
C139 x3.GN3 select2 0.00233f
C140 a_5699_5631# select0 9.55e-19
C141 x3.GN2 x5.GN 7.45e-19
C142 x3.GN2 x3.GN3 0.179278f
C143 VDD select0 1.13942f
C144 x5.A x5.GN 4.01022f
C145 x3.GN3 x5.A 0.430194f
C146 select2 x3.GN4 5.71e-20
C147 x3.GN2 x3.GN4 0.061048f
C148 x5.GN A1 0.558172f
C149 x3.GN3 A1 2.84e-19
C150 select2 select1 0.289185f
C151 a_5645_5493# select2 4.33e-19
C152 a_5645_7149# a_5699_7287# 0.006584f
C153 x5.GN x3.GP3 3.82e-20
C154 x3.GN3 x3.GP3 5.02512f
C155 x3.GN2 select1 0.108644f
C156 x5.A x3.GN4 0.446875f
C157 a_5645_5493# x3.GN2 0.039612f
C158 x3.GN4 A1 1.72e-19
C159 VDD A2 1.60691f
C160 A6 VDD 1.60651f
C161 x3.GN4 x3.GP3 5.65242f
C162 select1 A1 4.98e-22
C163 a_5699_5631# x3.GN1 0.001144f
C164 select1 x3.GP3 0.003325f
C165 a_5645_6637# x1.nSEL0 1.21e-20
C166 x3.GN1 VDD 0.890574f
C167 VDD a_5671_6589# 0.001496f
C168 x3.GN2 A7 0.006482f
C169 x4.A Z 5.48434f
C170 A6 A8 2.39e-19
C171 A7 x3.GP3 4.00999f
C172 a_5645_6637# a_5645_6461# 0.185422f
C173 a_5699_5631# VDD 9.09e-19
C174 x1.nSEL0 a_5645_6085# 0.001174f
C175 x1.nSEL1 select0 0.169954f
C176 A5 select2 2.94e-19
C177 A5 x3.GN2 0.145599f
C178 a_5645_6085# a_5645_5909# 0.185422f
C179 x1.nSEL0 a_5671_6037# 2.51e-19
C180 A5 x5.A 4.07e-21
C181 a_5645_5909# a_5671_6037# 0.004764f
C182 A5 x3.GP3 2.05e-19
C183 select2 select0 0.446748f
C184 x3.GN2 select0 0.114399f
C185 x4.A x5.GN 4.14756f
C186 x3.GN3 x4.A 0.430135f
C187 x3.GN1 x1.nSEL1 0.034871f
C188 VDD A8 1.54289f
C189 a_5645_6085# a_5645_6461# 3.02e-19
C190 x1.nSEL1 a_5671_6589# 4.08e-19
C191 select0 A1 2.25e-21
C192 x4.A x3.GN4 0.446815f
C193 x3.GP3 select0 2.74e-19
C194 x3.GN2 A2 3.77931f
C195 A6 x3.GN2 3.81318f
C196 x5.A A2 4.52052f
C197 x3.GN1 select2 0.054258f
C198 A1 A2 1.81909f
C199 x3.GN1 x3.GN2 0.146872f
C200 x3.GP3 A2 0.001569f
C201 x3.GN2 a_5671_6589# 3.11e-20
C202 A6 x3.GP3 0.001573f
C203 m2_5776_5494# x1.nSEL0 3.43e-19
C204 x3.GN3 A4 0.007342f
C205 x3.GN1 x5.A 0.43108f
C206 x3.GN1 A1 4.31229f
C207 a_5699_5631# x1.nSEL1 0.00175f
C208 x3.GN1 x3.GP3 0.076333f
C209 A4 x3.GN4 3.82686f
C210 VDD x1.nSEL1 0.472688f
C211 a_5671_6589# x3.GP3 4.39e-19
C212 x4.A A7 4.5214f
C213 a_5645_7149# x5.GN 1.19e-19
C214 x3.GN3 a_5645_7149# 1.07e-20
C215 a_5699_5631# x3.GN2 8.86e-19
C216 VDD select2 3.45811f
C217 VDD x3.GN2 0.700679f
C218 a_5645_7149# x3.GN4 0.134079f
C219 A3 x5.GN 7.03e-21
C220 A3 x3.GN3 3.78543f
C221 VDD x5.A 14.131701f
C222 a_5645_7149# select1 0.125445f
C223 VDD A1 1.63161f
C224 A5 x4.A 4.52088f
C225 A3 x3.GN4 0.16467f
C226 VDD x3.GP3 3.24607f
C227 x1.nSEL0 x5.GN 0.043717f
C228 x1.nSEL0 x3.GN3 4.01e-20
C229 x5.GN a_5645_5909# 3.56e-19
C230 x3.GN3 a_5645_5909# 6.68e-19
C231 x1.nSEL0 x3.GN4 2.26e-20
C232 x1.nSEL0 select1 0.137595f
C233 a_5645_5493# x1.nSEL0 0.081627f
C234 A5 A4 1.27332f
C235 select1 a_5645_5909# 0.03417f
C236 x3.GP3 A8 0.161339f
C237 a_5645_5493# a_5645_5909# 0.002207f
C238 A6 x4.A 4.52053f
C239 a_5645_6461# x5.GN 3.51e-19
C240 a_5645_6461# x3.GN3 0.104374f
C241 x3.GN1 x4.A 0.428411f
C242 a_5645_6461# x3.GN4 6.84e-19
C243 select2 x1.nSEL1 0.164995f
C244 x3.GN2 x1.nSEL1 0.209954f
C245 a_5645_6461# select1 0.261734f
C246 A4 A2 2.39e-19
C247 A6 A4 7.47e-20
C248 a_5645_7149# select0 0.220366f
C249 x3.GN2 select2 0.001516f
C250 x3.GN1 A4 0.218459f
C251 select2 x5.A 5.67943f
C252 x3.GN2 x5.A 0.429652f
C253 VDD x4.A 14.4067f
C254 select2 A1 0.054741f
C255 select2 x3.GP3 1.6e-19
C256 x3.GN2 A1 0.13437f
C257 x3.GN2 x3.GP3 0.060968f
C258 x5.A A1 4.52065f
C259 x5.A x3.GP3 0.358718f
C260 A3 A2 1.81997f
C261 x3.GP3 A1 1.96e-19
C262 x1.nSEL0 select0 0.325123f
C263 a_5645_6637# x5.GN 2.27e-19
C264 a_5645_6637# x3.GN3 0.004289f
C265 select0 a_5645_5909# 0.246189f
C266 Z VSS 6.934591f
C267 A8 VSS 3.687323f
C268 A7 VSS 3.163348f
C269 A6 VSS 3.279468f
C270 A5 VSS 3.50027f
C271 A4 VSS 3.017173f
C272 A3 VSS 3.199769f
C273 A2 VSS 4.079258f
C274 A1 VSS 5.727202f
C275 select2 VSS 6.977657f
C276 select0 VSS 1.45124f
C277 select1 VSS 1.80202f
C278 VDD VSS 0.118194p
C279 m2_5776_5494# VSS 0.065655f $ **FLOATING
C280 x4.A VSS 16.8199f
C281 x5.A VSS 13.867f
C282 a_5699_5631# VSS 0.006505f
C283 a_5645_5493# VSS 0.266782f
C284 x1.nSEL0 VSS 0.650696f
C285 x3.GN1 VSS 11.786012f
C286 a_5671_6037# VSS 0.004461f
C287 a_5645_5909# VSS 0.220868f
C288 x1.nSEL1 VSS 0.682637f
C289 x3.GN2 VSS 7.18136f
C290 a_5645_6085# VSS 0.23458f
C291 x5.GN VSS 5.83987f
C292 x3.GP3 VSS 3.19322f
C293 a_5671_6589# VSS 0.006801f
C294 x3.GN3 VSS 6.84829f
C295 a_5645_6461# VSS 0.232731f
C296 a_5645_6637# VSS 0.249604f
C297 x3.GN4 VSS 13.500038f
C298 a_5699_7287# VSS 0.006583f
C299 a_5645_7149# VSS 0.307391f
C300 x3.x2.GP VSS 3.41949f
C301 x2.x2.GP VSS 2.49707f
C302 x1.gpo1 VSS 0.984024f
C303 x3.GP2.t3 VSS 0.018013f
C304 x3.GP2.t2 VSS 0.018013f
C305 x3.GP2.n0 VSS 0.042951f
C306 x1.x12.Y VSS 0.065375f
C307 x3.GP2.n1 VSS 0.084381f
C308 x3.GP2.n2 VSS 0.026255f
C309 x3.GP2.t5 VSS 0.911601f
C310 x3.GP2.t7 VSS 0.937021f
C311 x3.GP2.n3 VSS 3.3244f
C312 x3.GP2.t4 VSS 0.911601f
C313 x3.GP2.t6 VSS 0.937021f
C314 x3.GP2.n4 VSS 3.3244f
C315 x3.GP2.n5 VSS 1.96615f
C316 x3.GP2.t1 VSS 0.027712f
C317 x3.GP2.t0 VSS 0.027712f
C318 x3.GP2.n6 VSS 0.057149f
C319 x3.GP2.n7 VSS 0.119653f
C320 A8.t1 VSS 0.893325f
C321 A8.t0 VSS 0.512841f
C322 A8.n0 VSS 4.96695f
C323 A8.t3 VSS 0.924602f
C324 A8.t2 VSS 0.65407f
C325 A8.n1 VSS 5.0783f
C326 A8.n2 VSS 0.803255f
C327 A8.n3 VSS 0.258761f
C328 A6.t2 VSS 0.763965f
C329 A6.t1 VSS 0.438578f
C330 A6.n0 VSS 4.2477f
C331 A6.t3 VSS 0.790712f
C332 A6.t0 VSS 0.559356f
C333 A6.n1 VSS 4.34292f
C334 A6.n2 VSS 0.686937f
C335 A6.n3 VSS 0.222065f
C336 A3.t1 VSS 0.893857f
C337 A3.t0 VSS 0.513146f
C338 A3.n0 VSS 4.9699f
C339 A3.t3 VSS 0.925152f
C340 A3.t2 VSS 0.654459f
C341 A3.n1 VSS 5.08132f
C342 A3.n2 VSS 0.803733f
C343 A3.n3 VSS 0.264783f
C344 A7.t1 VSS 0.893857f
C345 A7.t0 VSS 0.513146f
C346 A7.n0 VSS 4.9699f
C347 A7.t2 VSS 0.925152f
C348 A7.t3 VSS 0.654459f
C349 A7.n1 VSS 5.08132f
C350 A7.n2 VSS 0.803733f
C351 A7.n3 VSS 0.264783f
C352 A4.t1 VSS 0.893325f
C353 A4.t0 VSS 0.512841f
C354 A4.n0 VSS 4.96695f
C355 A4.t2 VSS 0.924602f
C356 A4.t3 VSS 0.65407f
C357 A4.n1 VSS 5.0783f
C358 A4.n2 VSS 0.803255f
C359 A4.n3 VSS 0.258761f
C360 A2.t1 VSS 0.763965f
C361 A2.t2 VSS 0.438578f
C362 A2.n0 VSS 4.2477f
C363 A2.t0 VSS 0.790712f
C364 A2.t3 VSS 0.559356f
C365 A2.n1 VSS 4.34292f
C366 A2.n2 VSS 0.686937f
C367 A2.n3 VSS 0.222065f
C368 A1.t2 VSS 0.795131f
C369 A1.t3 VSS 0.45647f
C370 A1.n0 VSS 4.42098f
C371 A1.t0 VSS 0.82297f
C372 A1.t1 VSS 0.582175f
C373 A1.n1 VSS 4.52009f
C374 A1.n2 VSS 0.714961f
C375 A1.n3 VSS 0.223162f
C376 x3.x1.GP VSS 3.39992f
C377 x2.GP1 VSS 2.31303f
C378 x1.gpo0 VSS 0.774629f
C379 x3.GP1.t3 VSS 0.01774f
C380 x3.GP1.t2 VSS 0.01774f
C381 x3.GP1.n0 VSS 0.0423f
C382 x1.x11.Y VSS 0.064713f
C383 x3.GP1.n1 VSS 0.083102f
C384 x3.GP1.n2 VSS 0.025857f
C385 x3.GP1.t6 VSS 0.897787f
C386 x3.GP1.t7 VSS 0.922822f
C387 x3.GP1.n3 VSS 3.26002f
C388 x3.GP1.t4 VSS 0.897787f
C389 x3.GP1.t5 VSS 0.922822f
C390 x3.GP1.n4 VSS 3.29215f
C391 x3.GP1.n5 VSS 1.7367f
C392 x3.GP1.t1 VSS 0.027292f
C393 x3.GP1.t0 VSS 0.027292f
C394 x3.GP1.n6 VSS 0.056236f
C395 x3.GP1.n7 VSS 0.120059f
C396 x3.x4.GP VSS 2.7871f
C397 x2.x4.GP VSS 2.18964f
C398 x1.gpo3 VSS 1.36452f
C399 x3.GP4.t2 VSS 0.01237f
C400 x3.GP4.t3 VSS 0.01237f
C401 x3.GP4.n0 VSS 0.029497f
C402 x1.x14.Y VSS 0.106916f
C403 x3.GP4.n1 VSS 0.056891f
C404 x3.GP4.t6 VSS 0.626043f
C405 x3.GP4.t4 VSS 0.643501f
C406 x3.GP4.n2 VSS 2.2877f
C407 x3.GP4.t5 VSS 0.626043f
C408 x3.GP4.t7 VSS 0.643501f
C409 x3.GP4.n3 VSS 2.2877f
C410 x3.GP4.n4 VSS 2.68712f
C411 x3.GP4.n5 VSS 0.0412f
C412 x3.GP4.n6 VSS 0.01803f
C413 x3.GP4.t0 VSS 0.019031f
C414 x3.GP4.t1 VSS 0.019031f
C415 x3.GP4.n7 VSS 0.041797f
C416 x3.GN4.t1 VSS 0.053314f
C417 x3.GN4.n0 VSS 0.061459f
C418 x3.GN4.t6 VSS 0.602506f
C419 x3.GN4.t9 VSS 0.587969f
C420 x3.GN4.n1 VSS 2.63799f
C421 x3.GN4.n2 VSS 1.63287f
C422 x3.GN4.t3 VSS 0.602506f
C423 x3.GN4.t5 VSS 0.587969f
C424 x3.GN4.n3 VSS 2.63799f
C425 x3.GN4.n4 VSS 2.31206f
C426 x3.GN4.t4 VSS 0.033468f
C427 x3.GN4.t2 VSS 0.019723f
C428 x3.GN4.t8 VSS 0.033468f
C429 x3.GN4.t7 VSS 0.019723f
C430 x3.GN4.n5 VSS 0.056155f
C431 x3.GN4.n6 VSS 0.083188f
C432 x3.GN4.n7 VSS 0.037242f
C433 x3.GN4.n8 VSS 0.301663f
C434 x3.GN4.t0 VSS 0.13616f
C435 x3.GN4.n9 VSS 0.024491f
C436 x3.GN4.n10 VSS 0.027436f
C437 A5.t2 VSS 0.770284f
C438 A5.t1 VSS 0.442205f
C439 A5.n0 VSS 4.28283f
C440 A5.t0 VSS 0.797252f
C441 A5.t3 VSS 0.563982f
C442 A5.n1 VSS 4.37884f
C443 A5.n2 VSS 0.692619f
C444 A5.n3 VSS 0.216188f
C445 x3.GN1.n0 VSS 1.21089f
C446 x3.GN1.t1 VSS 0.038044f
C447 x3.GN1.n1 VSS 0.0439f
C448 x3.GN1.t9 VSS 0.429934f
C449 x3.GN1.t7 VSS 0.419561f
C450 x3.GN1.n2 VSS 1.88241f
C451 x3.GN1.t2 VSS 0.429934f
C452 x3.GN1.t3 VSS 0.419561f
C453 x3.GN1.n3 VSS 1.88241f
C454 x3.GN1.n4 VSS 0.89272f
C455 x3.GN1.n5 VSS 0.303881f
C456 x3.GN1.t8 VSS 0.023882f
C457 x3.GN1.t5 VSS 0.014074f
C458 x3.GN1.t6 VSS 0.023882f
C459 x3.GN1.t4 VSS 0.014074f
C460 x3.GN1.n6 VSS 0.040071f
C461 x3.GN1.n7 VSS 0.059186f
C462 x3.GN1.n8 VSS 0.057565f
C463 x3.GN1.n9 VSS 0.125034f
C464 x3.GN1.t0 VSS 0.097161f
C465 x3.GN1.n10 VSS 0.017476f
C466 x3.GN1.n11 VSS 0.019578f
C467 VDD.n0 VSS 0.078152f
C468 VDD.n1 VSS 0.253693f
C469 VDD.n2 VSS 0.122926f
C470 VDD.n3 VSS 0.122926f
C471 VDD.n4 VSS 0.122525f
C472 VDD.n5 VSS 0.169863f
C473 VDD.n6 VSS 0.547624f
C474 VDD.t76 VSS 0.790353f
C475 VDD.n7 VSS 0.763087f
C476 VDD.t75 VSS 0.790353f
C477 VDD.n8 VSS 0.547624f
C478 VDD.n9 VSS 0.004814f
C479 VDD.n10 VSS 0.134493f
C480 VDD.n11 VSS 0.040318f
C481 VDD.n12 VSS 0.138067f
C482 VDD.n13 VSS 0.057005f
C483 VDD.n14 VSS 0.253704f
C484 VDD.n15 VSS 0.122531f
C485 VDD.n16 VSS 1.03197f
C486 VDD.n17 VSS 1.03197f
C487 VDD.n18 VSS 0.169845f
C488 VDD.n19 VSS 0.124397f
C489 VDD.t22 VSS 1.37216f
C490 VDD.n22 VSS 0.124397f
C491 VDD.n23 VSS 5.27e-19
C492 VDD.n24 VSS 0.07554f
C493 VDD.n25 VSS 0.013735f
C494 VDD.n26 VSS 0.149327f
C495 VDD.n27 VSS 0.079843f
C496 VDD.n28 VSS 0.162134f
C497 VDD.n29 VSS 0.188097f
C498 VDD.n30 VSS 0.253704f
C499 VDD.n31 VSS 0.004119f
C500 VDD.n32 VSS 0.169845f
C501 VDD.n33 VSS 0.124397f
C502 VDD.t41 VSS 1.37216f
C503 VDD.n35 VSS 1.03197f
C504 VDD.n36 VSS 0.124397f
C505 VDD.n38 VSS 1.03197f
C506 VDD.n39 VSS 0.122531f
C507 VDD.n40 VSS 0.009862f
C508 VDD.n41 VSS 0.075465f
C509 VDD.n42 VSS 0.013861f
C510 VDD.n43 VSS 0.149327f
C511 VDD.n44 VSS 0.079211f
C512 VDD.n45 VSS 0.128376f
C513 VDD.n46 VSS 0.184404f
C514 VDD.n47 VSS 0.253704f
C515 VDD.n48 VSS 0.00437f
C516 VDD.n49 VSS 0.169845f
C517 VDD.n50 VSS 0.124397f
C518 VDD.t7 VSS 1.37216f
C519 VDD.n52 VSS 1.03197f
C520 VDD.n53 VSS 0.124397f
C521 VDD.n55 VSS 1.03197f
C522 VDD.n56 VSS 0.122531f
C523 VDD.n57 VSS 0.009878f
C524 VDD.n58 VSS 0.075214f
C525 VDD.n59 VSS 0.013861f
C526 VDD.n60 VSS 0.149327f
C527 VDD.n61 VSS 0.079211f
C528 VDD.n62 VSS 0.125941f
C529 VDD.n63 VSS 0.167914f
C530 VDD.n64 VSS 0.010164f
C531 VDD.n65 VSS 0.00773f
C532 VDD.t32 VSS 0.015599f
C533 VDD.n66 VSS 0.015344f
C534 VDD.t52 VSS 0.001675f
C535 VDD.t21 VSS 0.002544f
C536 VDD.n67 VSS 0.004395f
C537 VDD.t30 VSS 0.015899f
C538 VDD.t74 VSS 0.015599f
C539 VDD.n68 VSS 0.014858f
C540 VDD.n69 VSS 0.00773f
C541 VDD.n70 VSS 0.006997f
C542 VDD.t9 VSS 0.002296f
C543 VDD.n71 VSS 0.006515f
C544 VDD.t60 VSS 0.009437f
C545 VDD.n72 VSS 0.008687f
C546 VDD.n73 VSS 0.007753f
C547 VDD.t26 VSS 0.015603f
C548 VDD.n74 VSS 0.001276f
C549 VDD.t47 VSS 0.00669f
C550 VDD.t62 VSS 0.011043f
C551 VDD.n75 VSS 0.010887f
C552 VDD.n76 VSS 0.013048f
C553 VDD.t79 VSS 0.046088f
C554 VDD.n77 VSS 0.041686f
C555 VDD.t38 VSS 0.00125f
C556 VDD.t44 VSS 0.003352f
C557 VDD.n78 VSS 0.0153f
C558 VDD.t63 VSS 0.011043f
C559 VDD.n79 VSS 0.008081f
C560 VDD.n80 VSS 0.030158f
C561 VDD.n81 VSS 0.023827f
C562 VDD.n82 VSS 0.030949f
C563 VDD.n83 VSS 0.01787f
C564 VDD.n84 VSS 0.013048f
C565 VDD.n85 VSS 0.009786f
C566 VDD.n86 VSS 0.006143f
C567 VDD.n87 VSS 0.019352f
C568 VDD.n88 VSS 0.030339f
C569 VDD.t39 VSS 0.031357f
C570 VDD.n89 VSS 0.002361f
C571 VDD.n90 VSS 0.002411f
C572 VDD.n91 VSS 0.009786f
C573 VDD.n92 VSS 0.003014f
C574 VDD.t24 VSS 0.015814f
C575 VDD.n93 VSS 0.012977f
C576 VDD.n94 VSS 0.00773f
C577 VDD.t80 VSS 0.046088f
C578 VDD.n95 VSS 0.011488f
C579 VDD.n96 VSS 0.00773f
C580 VDD.t36 VSS 0.00125f
C581 VDD.t49 VSS 0.003352f
C582 VDD.n97 VSS 0.0153f
C583 VDD.t82 VSS 0.046088f
C584 VDD.t56 VSS 0.00669f
C585 VDD.n98 VSS 0.020658f
C586 VDD.n99 VSS 0.011843f
C587 VDD.n100 VSS 0.006143f
C588 VDD.t65 VSS 0.011043f
C589 VDD.n101 VSS 0.010887f
C590 VDD.n102 VSS 0.041686f
C591 VDD.n103 VSS 0.01787f
C592 VDD.n104 VSS 0.030949f
C593 VDD.t66 VSS 0.011043f
C594 VDD.t34 VSS 0.015815f
C595 VDD.n105 VSS 0.004468f
C596 VDD.n106 VSS 0.005319f
C597 VDD.t55 VSS 0.063133f
C598 VDD.t48 VSS 0.061042f
C599 VDD.t64 VSS 0.045154f
C600 VDD.t35 VSS 0.064805f
C601 VDD.t11 VSS 0.063133f
C602 VDD.t13 VSS 0.071913f
C603 VDD.t15 VSS 0.052262f
C604 VDD.t27 VSS 0.028013f
C605 VDD.t23 VSS 0.012961f
C606 VDD.t33 VSS 0.045572f
C607 VDD.n107 VSS 0.059469f
C608 VDD.n108 VSS 0.041241f
C609 VDD.n109 VSS 0.012122f
C610 VDD.n110 VSS 0.01945f
C611 VDD.n111 VSS 0.023827f
C612 VDD.n112 VSS 0.008084f
C613 VDD.n113 VSS 0.064395f
C614 VDD.n114 VSS 0.087594f
C615 VDD.t71 VSS 0.011043f
C616 VDD.n115 VSS 0.021596f
C617 VDD.n116 VSS 0.041686f
C618 VDD.n117 VSS 0.025689f
C619 VDD.t72 VSS 0.011043f
C620 VDD.t1 VSS 0.015891f
C621 VDD.n118 VSS 0.018568f
C622 VDD.t70 VSS 0.142033f
C623 VDD.t67 VSS 0.087258f
C624 VDD.t18 VSS 0.035804f
C625 VDD.t77 VSS 0.049557f
C626 VDD.t53 VSS 0.035804f
C627 VDD.t57 VSS 0.049557f
C628 VDD.t3 VSS 0.035804f
C629 VDD.t0 VSS 0.053589f
C630 VDD.n119 VSS 0.058661f
C631 VDD.n120 VSS 0.00773f
C632 VDD.n121 VSS 0.003365f
C633 VDD.t58 VSS 0.015891f
C634 VDD.n122 VSS 0.003365f
C635 VDD.t78 VSS 0.015891f
C636 VDD.n123 VSS 0.227132f
C637 VDD.n124 VSS 0.013294f
C638 VDD.n125 VSS 0.008081f
C639 VDD.t81 VSS 0.046809f
C640 VDD.t68 VSS 0.011043f
C641 VDD.n126 VSS 0.04634f
C642 VDD.n127 VSS 0.023029f
C643 VDD.t69 VSS 0.011043f
C644 VDD.n128 VSS 0.030158f
C645 VDD.n129 VSS 0.027736f
C646 VDD.n130 VSS 0.017403f
C647 VDD.n131 VSS 0.013581f
C648 VDD.n132 VSS 0.013243f
C649 VDD.t19 VSS 0.015899f
C650 VDD.n133 VSS 0.020008f
C651 VDD.n134 VSS 0.00773f
C652 VDD.n135 VSS 0.013048f
C653 VDD.n136 VSS 0.009786f
C654 VDD.n137 VSS 0.018769f
C655 VDD.t54 VSS 0.015899f
C656 VDD.n138 VSS 0.02031f
C657 VDD.n139 VSS 0.00773f
C658 VDD.n140 VSS 0.013048f
C659 VDD.n141 VSS 0.009786f
C660 VDD.n142 VSS 0.018769f
C661 VDD.t4 VSS 0.015899f
C662 VDD.n143 VSS 0.02031f
C663 VDD.n144 VSS 0.003365f
C664 VDD.n145 VSS 0.013048f
C665 VDD.n146 VSS 0.009786f
C666 VDD.n147 VSS 0.004964f
C667 VDD.n148 VSS 0.027117f
C668 VDD.n149 VSS 0.012122f
C669 VDD.n150 VSS 0.01945f
C670 VDD.n151 VSS 0.033134f
C671 VDD.n152 VSS 0.006595f
C672 VDD.n153 VSS 0.059927f
C673 VDD.n154 VSS 0.058109f
C674 VDD.n155 VSS 0.001347f
C675 VDD.t28 VSS 0.001675f
C676 VDD.t16 VSS 0.002544f
C677 VDD.n156 VSS 0.004395f
C678 VDD.n157 VSS 0.029498f
C679 VDD.t14 VSS 0.015891f
C680 VDD.n158 VSS 0.018518f
C681 VDD.t50 VSS 0.005236f
C682 VDD.t40 VSS 0.013917f
C683 VDD.n159 VSS 0.007895f
C684 VDD.t12 VSS 0.015603f
C685 VDD.n160 VSS 0.016462f
C686 VDD.n161 VSS 0.021174f
C687 VDD.n162 VSS 0.002788f
C688 VDD.n163 VSS 0.013048f
C689 VDD.n164 VSS 0.00773f
C690 VDD.n165 VSS 0.004468f
C691 VDD.n166 VSS 0.004964f
C692 VDD.n167 VSS 0.026569f
C693 VDD.n168 VSS 0.072449f
C694 VDD.t51 VSS 0.013797f
C695 VDD.t31 VSS 0.035956f
C696 VDD.t29 VSS 0.040137f
C697 VDD.t20 VSS 0.028013f
C698 VDD.t8 VSS 0.052262f
C699 VDD.t73 VSS 0.073585f
C700 VDD.t25 VSS 0.035956f
C701 VDD.t59 VSS 0.028013f
C702 VDD.t37 VSS 0.064805f
C703 VDD.t61 VSS 0.045154f
C704 VDD.t43 VSS 0.061042f
C705 VDD.t46 VSS 0.063133f
C706 VDD.n169 VSS 0.042993f
C707 VDD.n170 VSS 0.01249f
C708 VDD.n171 VSS 0.008891f
C709 VDD.n172 VSS 0.002361f
C710 VDD.n173 VSS 0.017322f
C711 VDD.n174 VSS 0.006606f
C712 VDD.n175 VSS 0.013048f
C713 VDD.n176 VSS 0.009786f
C714 VDD.n177 VSS 0.005817f
C715 VDD.n178 VSS 0.019774f
C716 VDD.n179 VSS 0.014151f
C717 VDD.n180 VSS 0.009006f
C718 VDD.n181 VSS 0.025467f
C719 VDD.n182 VSS 0.279991f
C720 VDD.n183 VSS 0.651519f
C721 VDD.n184 VSS 0.253704f
C722 VDD.n185 VSS 0.051921f
C723 VDD.n186 VSS 0.122531f
C724 VDD.n187 VSS 1.03197f
C725 VDD.n188 VSS 1.03197f
C726 VDD.n189 VSS 0.169845f
C727 VDD.n190 VSS 0.124397f
C728 VDD.t45 VSS 1.37216f
C729 VDD.n193 VSS 0.124397f
C730 VDD.n194 VSS 4.77e-19
C731 VDD.n195 VSS 0.07554f
C732 VDD.n196 VSS 0.013785f
C733 VDD.n197 VSS 0.149327f
C734 VDD.n198 VSS 0.079793f
C735 VDD.n199 VSS 0.15219f
C736 VDD.n200 VSS 0.253704f
C737 VDD.n201 VSS 0.00437f
C738 VDD.n202 VSS 0.169845f
C739 VDD.n203 VSS 0.124397f
C740 VDD.t17 VSS 1.37216f
C741 VDD.n205 VSS 1.03197f
C742 VDD.n206 VSS 0.124397f
C743 VDD.n208 VSS 1.03197f
C744 VDD.n209 VSS 0.122531f
C745 VDD.n210 VSS 0.075214f
C746 VDD.n211 VSS 0.013861f
C747 VDD.n212 VSS 0.149327f
C748 VDD.n213 VSS 0.079211f
C749 VDD.n214 VSS 0.153404f
C750 VDD.n215 VSS 0.196603f
C751 VDD.n216 VSS 0.116414f
C752 VDD.n217 VSS 0.075465f
C753 VDD.n218 VSS 0.013861f
C754 VDD.n219 VSS 1.03197f
C755 VDD.n220 VSS 1.03197f
C756 VDD.n221 VSS 0.122531f
C757 VDD.n222 VSS 0.079211f
C758 VDD.n223 VSS 0.149327f
C759 VDD.n224 VSS 0.253704f
C760 VDD.n225 VSS 0.169845f
C761 VDD.n226 VSS 0.124397f
C762 VDD.t42 VSS 1.37216f
C763 VDD.n229 VSS 0.124397f
C764 VDD.n230 VSS 0.004119f
C765 VDD.n231 VSS 0.009862f
C766 VDD.n232 VSS 0.235683f
C767 VDD.n233 VSS 0.097082f
C768 VDD.n234 VSS 5.27e-19
C769 VDD.n235 VSS 0.079843f
C770 VDD.n236 VSS 0.149327f
C771 VDD.n237 VSS 0.169845f
C772 VDD.n238 VSS 0.124397f
C773 VDD.t10 VSS 1.37216f
C774 VDD.n239 VSS 0.253704f
C775 VDD.n241 VSS 1.03197f
C776 VDD.n242 VSS 0.124397f
C777 VDD.n244 VSS 1.03197f
C778 VDD.n245 VSS 0.122531f
C779 VDD.n246 VSS 0.07554f
C780 VDD.n247 VSS 0.013735f
C781 VDD.n248 VSS 0.013528f
C782 VDD.n249 VSS 0.191035f
C783 VDD.n250 VSS 0.253704f
C784 VDD.n251 VSS 0.07554f
C785 VDD.n252 VSS 1.03197f
C786 VDD.n253 VSS 1.03197f
C787 VDD.n254 VSS 0.122531f
C788 VDD.n255 VSS 0.169845f
C789 VDD.n256 VSS 0.124397f
C790 VDD.t6 VSS 1.37216f
C791 VDD.n259 VSS 0.124397f
C792 VDD.n260 VSS 4.77e-19
C793 VDD.n261 VSS 0.013492f
C794 VDD.n262 VSS 0.013785f
C795 VDD.n263 VSS 0.149327f
C796 VDD.n264 VSS 0.079793f
C797 VDD.n265 VSS 0.142932f
C798 VDD.n266 VSS 0.154755f
C799 VDD.n267 VSS 0.390936f
C800 VDD.n268 VSS 0.078152f
C801 VDD.n269 VSS 0.253693f
C802 VDD.n270 VSS 0.122926f
C803 VDD.n271 VSS 0.122926f
C804 VDD.n272 VSS 0.122525f
C805 VDD.n273 VSS 0.169863f
C806 VDD.n274 VSS 0.547624f
C807 VDD.t2 VSS 0.790353f
C808 VDD.n275 VSS 0.763087f
C809 VDD.t5 VSS 0.790353f
C810 VDD.n276 VSS 0.547624f
C811 VDD.n277 VSS 0.004814f
C812 VDD.n278 VSS 0.134493f
C813 VDD.n279 VSS 0.040288f
C814 VDD.n280 VSS 0.072753f
C815 Z.t1 VSS 0.434416f
C816 Z.n0 VSS 0.540283f
C817 Z.t0 VSS 0.446377f
C818 Z.t5 VSS 0.336375f
C819 Z.n1 VSS 2.25255f
C820 Z.n2 VSS 0.762169f
C821 Z.t4 VSS 0.329756f
C822 Z.n3 VSS 0.492384f
C823 Z.n4 VSS 0.648657f
C824 Z.n5 VSS 0.805956f
C825 Z.t6 VSS 0.434416f
C826 Z.n6 VSS 0.540283f
C827 Z.t7 VSS 0.446377f
C828 Z.t2 VSS 0.336375f
C829 Z.n7 VSS 2.25255f
C830 Z.n8 VSS 0.762169f
C831 Z.t3 VSS 0.329756f
C832 Z.n9 VSS 0.492384f
C833 Z.n10 VSS 0.664311f
C834 Z.n11 VSS 0.690962f
C835 select2.t3 VSS 0.587177f
C836 select2.t4 VSS 0.57301f
C837 select2.n0 VSS 2.59538f
C838 select2.t1 VSS 0.032617f
C839 select2.t7 VSS 0.019221f
C840 select2.t6 VSS 0.032617f
C841 select2.t5 VSS 0.019221f
C842 select2.n1 VSS 0.054727f
C843 select2.n2 VSS 0.080908f
C844 select2.n3 VSS 0.080265f
C845 select2.n4 VSS 1.30544f
C846 select2.t2 VSS 0.689751f
C847 select2.t0 VSS 0.708986f
C848 select2.n5 VSS 2.58319f
C849 select2.n6 VSS 1.73421f
C850 select2.n7 VSS 4.54326f
C851 select2.n8 VSS 1.57054f
C852 select1.t6 VSS 0.031316f
C853 select1.t5 VSS 0.018454f
C854 select1.t3 VSS 0.031316f
C855 select1.t1 VSS 0.018454f
C856 select1.n0 VSS 0.052544f
C857 select1.n1 VSS 0.077632f
C858 select1.n2 VSS 0.047269f
C859 select1.t9 VSS 0.014491f
C860 select1.t7 VSS 0.03056f
C861 select1.n3 VSS 0.109737f
C862 select1.n4 VSS 0.021277f
C863 select1.n5 VSS 0.018327f
C864 select1.t4 VSS 0.022078f
C865 select1.t2 VSS 0.015172f
C866 select1.n6 VSS 0.064155f
C867 select1.n7 VSS 0.014778f
C868 select1.n8 VSS 0.105859f
C869 select1.n9 VSS 0.383423f
C870 select1.t8 VSS 0.026898f
C871 select1.t0 VSS 0.018264f
C872 select1.n10 VSS 0.063549f
C873 select1.n11 VSS 0.015211f
C874 select1.n12 VSS 0.098666f
C875 select1.n13 VSS 0.442567f
C876 select1.n14 VSS 0.578172f
.ends

